//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1318, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G97), .C2(G257), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G1), .B2(G20), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n207), .B(new_n220), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT65), .B(G250), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n231), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G116), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT69), .B(G107), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n221), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT72), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n255), .A3(new_n221), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n204), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n257), .A2(G50), .A3(new_n249), .A4(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G58), .ZN(new_n262));
  INV_X1    g0062(.A(G58), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT8), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT73), .ZN(new_n265));
  OR3_X1    g0065(.A1(new_n263), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n204), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G150), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n269), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT74), .B1(new_n269), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G58), .A2(G68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n204), .B1(new_n274), .B2(new_n213), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n251), .B(new_n260), .C1(new_n276), .C2(new_n257), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT71), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n279), .A2(new_n281), .A3(new_n284), .A4(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(G223), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n279), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G77), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n289), .A2(new_n293), .A3(G222), .A4(new_n290), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n286), .A2(new_n288), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n203), .B(G274), .C1(G41), .C2(G45), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n214), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n277), .B1(G179), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n277), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n260), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n269), .A2(new_n271), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n275), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n269), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n257), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT9), .A3(new_n251), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n305), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(new_n300), .ZN(new_n322));
  AOI211_X1 g0122(.A(new_n322), .B(new_n303), .C1(new_n295), .C2(new_n298), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G190), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n310), .A2(new_n320), .A3(new_n321), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n250), .B(new_n311), .C1(new_n317), .C2(new_n318), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(KEYINPUT9), .B1(G190), .B2(new_n323), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT10), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n321), .A4(new_n310), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n308), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n270), .A2(G50), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n215), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n267), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n336));
  NAND3_X1  g0136(.A1(new_n318), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n254), .A3(new_n256), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n203), .A2(new_n215), .A3(G13), .A4(G20), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g0145(.A(new_n249), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n253), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n249), .A2(KEYINPUT76), .A3(new_n221), .A4(new_n252), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n215), .B(new_n258), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n297), .A2(G238), .A3(new_n301), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G232), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G1698), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n289), .B1(G33), .B2(G97), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n300), .B(new_n353), .C1(new_n357), .C2(new_n297), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n214), .A2(new_n290), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(G1698), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n279), .A2(new_n360), .A3(new_n281), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n322), .B1(new_n364), .B2(new_n298), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n353), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n359), .A2(G179), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n359), .A2(new_n367), .A3(KEYINPUT79), .A4(G179), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n365), .B2(new_n353), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n297), .B1(new_n362), .B2(new_n363), .ZN(new_n374));
  INV_X1    g0174(.A(new_n353), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT13), .A4(new_n322), .ZN(new_n376));
  OAI21_X1  g0176(.A(G169), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n359), .A2(new_n367), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT14), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n372), .A2(new_n382), .A3(KEYINPUT80), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n379), .B2(G169), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT14), .B(new_n307), .C1(new_n359), .C2(new_n367), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n370), .A2(new_n371), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n352), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n379), .A2(G200), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n351), .C1(new_n392), .C2(new_n379), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n283), .A2(G238), .A3(new_n285), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n287), .A2(G107), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n298), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n297), .A2(G244), .A3(new_n301), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n300), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n322), .B1(new_n397), .B2(new_n298), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(G200), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT8), .B(G58), .ZN(new_n406));
  INV_X1    g0206(.A(new_n270), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT15), .B(G87), .Z(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n406), .A2(new_n407), .B1(new_n409), .B2(new_n267), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n204), .A2(new_n334), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n253), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n346), .A2(new_n334), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n347), .A2(new_n348), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(G77), .A3(new_n259), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n405), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT77), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n392), .B1(new_n402), .B2(new_n404), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n417), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n331), .A2(new_n390), .A3(new_n393), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n300), .B1(new_n302), .B2(new_n355), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT83), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n214), .A2(G1698), .ZN(new_n428));
  OR2_X1    g0228(.A1(G223), .A2(G1698), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n279), .A4(new_n281), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n298), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT83), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n300), .C1(new_n302), .C2(new_n355), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n427), .A2(new_n433), .A3(new_n392), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT84), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n297), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n426), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n436), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n265), .A2(new_n266), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n257), .B2(new_n249), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n263), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n406), .B2(KEYINPUT73), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n346), .B1(new_n447), .B2(new_n259), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT82), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n256), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n255), .B1(new_n252), .B2(new_n221), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n249), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n249), .B1(new_n444), .B2(new_n258), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(G58), .B(G68), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(G20), .B1(G159), .B2(new_n270), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n280), .A2(G33), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n204), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT7), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G20), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n462), .A2(new_n463), .B1(new_n287), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT16), .B(new_n459), .C1(new_n465), .C2(new_n215), .ZN(new_n466));
  INV_X1    g0266(.A(new_n459), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n280), .A2(KEYINPUT81), .A3(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n279), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n463), .B1(new_n289), .B2(G20), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n467), .B1(new_n474), .B2(G68), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n466), .B(new_n253), .C1(new_n475), .C2(KEYINPUT16), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n457), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT85), .B1(new_n443), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n436), .A2(new_n440), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT84), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n449), .A2(new_n456), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n475), .A2(KEYINPUT16), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n466), .A2(new_n253), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT85), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n478), .A2(new_n488), .A3(KEYINPUT17), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT18), .ZN(new_n490));
  INV_X1    g0290(.A(G179), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n427), .A2(new_n433), .A3(new_n491), .A4(new_n435), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n307), .B1(new_n439), .B2(new_n426), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n477), .A2(KEYINPUT18), .A3(new_n493), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n482), .A2(new_n486), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT17), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n489), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT75), .B1(new_n403), .B2(new_n399), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n491), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n402), .A2(new_n307), .A3(new_n404), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n416), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n425), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G303), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n287), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n290), .A2(G257), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G264), .A2(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n279), .A2(new_n281), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n298), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n203), .A2(G45), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G274), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n203), .B(G45), .C1(new_n522), .C2(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G270), .A3(new_n297), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G169), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n203), .A2(G33), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT91), .B1(new_n414), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT91), .ZN(new_n532));
  AOI211_X1 g0332(.A(new_n532), .B(new_n529), .C1(new_n347), .C2(new_n348), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n204), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT86), .B(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n278), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n209), .A2(G20), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n253), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n537), .ZN(new_n543));
  INV_X1    g0343(.A(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n548), .B2(G33), .ZN(new_n549));
  INV_X1    g0349(.A(new_n541), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT20), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n346), .A2(new_n209), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n527), .B1(new_n534), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n552), .B(new_n553), .C1(new_n531), .C2(new_n533), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n527), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n252), .A2(new_n221), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT76), .B1(new_n560), .B2(new_n249), .ZN(new_n561));
  INV_X1    g0361(.A(new_n348), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n530), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n532), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n414), .A2(KEYINPUT91), .A3(new_n530), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n542), .A2(new_n551), .B1(new_n209), .B2(new_n346), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n525), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n556), .A2(new_n559), .B1(G179), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n279), .B(new_n281), .C1(G250), .C2(G1698), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n290), .A2(G257), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT95), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT95), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n576), .A3(new_n298), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n523), .A2(new_n297), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G264), .B1(G274), .B2(new_n520), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n580), .A3(G179), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G107), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n585), .A2(KEYINPUT23), .A3(G20), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT23), .B1(new_n585), .B2(G20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n586), .A2(new_n587), .B1(G20), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT92), .A2(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n289), .A2(new_n204), .A3(G87), .A4(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n279), .A2(new_n281), .A3(new_n204), .A4(G87), .ZN(new_n592));
  INV_X1    g0392(.A(new_n590), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI211_X1 g0394(.A(KEYINPUT24), .B(new_n589), .C1(new_n591), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n591), .ZN(new_n597));
  INV_X1    g0397(.A(new_n589), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n253), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n346), .A2(new_n585), .ZN(new_n603));
  NOR2_X1   g0403(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n346), .A2(KEYINPUT93), .A3(KEYINPUT25), .A4(new_n585), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n257), .A2(new_n249), .A3(new_n528), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n585), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n600), .A2(new_n601), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n601), .B1(new_n600), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n584), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n581), .A2(G200), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n577), .A2(new_n580), .A3(G190), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n600), .A3(new_n610), .A4(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n557), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n525), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n618), .C1(new_n392), .C2(new_n525), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n569), .A2(new_n613), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n279), .A2(new_n281), .A3(G244), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT4), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n624), .A3(new_n536), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n289), .A2(G250), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n290), .B1(new_n626), .B2(KEYINPUT4), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n298), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n521), .B1(new_n578), .B2(new_n227), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n438), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n630), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n631), .A2(KEYINPUT88), .B1(new_n632), .B2(new_n392), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n249), .A2(G97), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n608), .B2(new_n544), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n463), .A2(new_n462), .B1(new_n471), .B2(new_n464), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n585), .ZN(new_n639));
  XOR2_X1   g0439(.A(G97), .B(G107), .Z(new_n640));
  NAND2_X1  g0440(.A1(new_n585), .A2(KEYINPUT6), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n640), .A2(KEYINPUT6), .B1(new_n548), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(G20), .B1(G77), .B2(new_n270), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n474), .A2(KEYINPUT87), .A3(G107), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n636), .B1(new_n645), .B2(new_n253), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n622), .A2(new_n623), .B1(G33), .B2(G283), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n623), .B1(new_n289), .B2(G250), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n647), .B(new_n621), .C1(new_n290), .C2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n629), .B1(new_n649), .B2(new_n298), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT88), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(G190), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n633), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n253), .ZN(new_n654));
  INV_X1    g0454(.A(new_n636), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n628), .A2(new_n491), .A3(new_n630), .ZN(new_n657));
  AOI21_X1  g0457(.A(G169), .B1(new_n628), .B2(new_n630), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n408), .A2(new_n249), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n289), .A2(new_n204), .A3(G68), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT19), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n548), .B2(new_n267), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n538), .A2(G87), .A3(G107), .ZN(new_n665));
  NAND3_X1  g0465(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n204), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n662), .B(new_n664), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n661), .B1(new_n668), .B2(new_n253), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n216), .A2(new_n290), .ZN(new_n670));
  INV_X1    g0470(.A(G244), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G1698), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n279), .A2(new_n670), .A3(new_n281), .A4(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n297), .B1(new_n673), .B2(new_n588), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n297), .A2(G250), .A3(new_n516), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n203), .A2(G45), .A3(G274), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G190), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(G238), .A2(G1698), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n671), .B2(G1698), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(new_n289), .B1(G33), .B2(G116), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n678), .B(new_n675), .C1(new_n682), .C2(new_n297), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G200), .ZN(new_n684));
  INV_X1    g0484(.A(new_n608), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G87), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n669), .A2(new_n679), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(G169), .ZN(new_n688));
  INV_X1    g0488(.A(new_n674), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(G179), .A3(new_n678), .A4(new_n675), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT89), .ZN(new_n692));
  INV_X1    g0492(.A(new_n661), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n257), .A2(new_n249), .A3(new_n408), .A4(new_n528), .ZN(new_n694));
  AOI21_X1  g0494(.A(G87), .B1(new_n545), .B2(new_n547), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n667), .B1(new_n695), .B2(new_n585), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n287), .A2(G20), .A3(new_n215), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT19), .B1(new_n538), .B2(new_n268), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n693), .B(new_n694), .C1(new_n699), .C2(new_n560), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n669), .A2(KEYINPUT90), .A3(new_n694), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n688), .A2(new_n704), .A3(new_n690), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n692), .A2(new_n702), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n653), .A2(new_n660), .A3(new_n687), .A4(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n509), .A2(new_n620), .A3(new_n707), .ZN(G372));
  AND4_X1   g0508(.A1(new_n504), .A2(new_n393), .A3(new_n505), .A4(new_n416), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT80), .B1(new_n372), .B2(new_n382), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n387), .A2(new_n384), .A3(new_n388), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n352), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n489), .A2(new_n500), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n497), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n326), .A2(new_n330), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n308), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n691), .A2(new_n700), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n687), .ZN(new_n720));
  AND4_X1   g0520(.A1(new_n616), .A2(new_n653), .A3(new_n660), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n597), .A2(new_n598), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT24), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n597), .A2(new_n596), .A3(new_n598), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n560), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n584), .B1(new_n725), .B2(new_n609), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n569), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n719), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(new_n687), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n628), .A2(new_n491), .A3(new_n630), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n650), .B2(G169), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n729), .A2(new_n646), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT96), .B1(new_n732), .B2(KEYINPUT26), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n646), .A2(new_n731), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n706), .A3(KEYINPUT26), .A4(new_n687), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n656), .A2(new_n659), .A3(new_n687), .A4(new_n718), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT26), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n717), .B1(new_n742), .B2(new_n509), .ZN(G369));
  OAI21_X1  g0543(.A(KEYINPUT94), .B1(new_n725), .B2(new_n609), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n600), .A2(new_n601), .A3(new_n610), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(new_n582), .B2(new_n583), .ZN(new_n746));
  INV_X1    g0546(.A(G13), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n203), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT27), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT27), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G213), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G343), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n613), .A2(new_n616), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n756), .B1(new_n611), .B2(new_n612), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n569), .A2(new_n756), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n756), .A2(new_n726), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n568), .A2(G179), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n558), .B1(new_n557), .B2(new_n527), .ZN(new_n769));
  AOI211_X1 g0569(.A(KEYINPUT21), .B(new_n526), .C1(new_n566), .C2(new_n567), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n619), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n617), .B2(new_n755), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n768), .B1(new_n770), .B2(new_n769), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n557), .A3(new_n756), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n762), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n779), .ZN(G399));
  NAND2_X1  g0580(.A1(new_n665), .A2(new_n209), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n205), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G41), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(G1), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n223), .B2(new_n785), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  INV_X1    g0588(.A(G330), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT30), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n683), .A2(new_n491), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(new_n580), .A3(new_n577), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n628), .A2(new_n524), .A3(new_n630), .A4(new_n515), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n795));
  OR3_X1    g0595(.A1(new_n792), .A2(new_n790), .A3(new_n793), .ZN(new_n796));
  AOI21_X1  g0596(.A(G179), .B1(new_n677), .B2(new_n678), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n581), .A2(new_n632), .A3(new_n797), .A4(new_n525), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT99), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(KEYINPUT31), .B1(new_n801), .B2(new_n756), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n620), .A2(new_n707), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n755), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n796), .A2(new_n798), .A3(new_n794), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(KEYINPUT31), .A3(new_n756), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n789), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT29), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n734), .A2(new_n706), .A3(new_n738), .A4(new_n687), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n719), .B1(new_n736), .B2(KEYINPUT26), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n746), .A2(new_n774), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n653), .A2(new_n660), .A3(new_n616), .A4(new_n720), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n809), .B1(new_n814), .B2(new_n755), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n756), .B1(new_n728), .B2(new_n740), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n788), .B1(new_n819), .B2(G1), .ZN(G364));
  NAND2_X1  g0620(.A1(new_n748), .A2(G45), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n785), .A2(G1), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n777), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n776), .A2(G330), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n221), .B1(G20), .B2(new_n307), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n204), .A2(G179), .ZN(new_n827));
  NOR2_X1   g0627(.A1(G190), .A2(G200), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n204), .A2(new_n491), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n835), .A3(new_n828), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n392), .A2(G200), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n834), .A2(new_n837), .A3(new_n835), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n832), .B1(new_n334), .B2(new_n836), .C1(new_n839), .C2(new_n263), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n491), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G20), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n544), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n833), .A2(G200), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(G190), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(G68), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n827), .A2(G190), .A3(G200), .ZN(new_n850));
  INV_X1    g0650(.A(G87), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n827), .A2(new_n392), .A3(G200), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n287), .B(new_n852), .C1(G107), .C2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n848), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n845), .A2(new_n392), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n840), .B(new_n856), .C1(G50), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n289), .B1(new_n842), .B2(G294), .ZN(new_n859));
  INV_X1    g0659(.A(G311), .ZN(new_n860));
  INV_X1    g0660(.A(G322), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n859), .B1(new_n860), .B2(new_n836), .C1(new_n839), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n850), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n857), .A2(G326), .B1(new_n865), .B2(G303), .ZN(new_n866));
  INV_X1    g0666(.A(G317), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT33), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(KEYINPUT33), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n846), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n829), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n872), .A2(G329), .ZN(new_n873));
  NOR4_X1   g0673(.A1(new_n862), .A2(new_n864), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n826), .B1(new_n858), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n783), .A2(new_n289), .ZN(new_n876));
  INV_X1    g0676(.A(G45), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n224), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n876), .B(new_n878), .C1(new_n243), .C2(new_n877), .ZN(new_n879));
  INV_X1    g0679(.A(G355), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n289), .A2(new_n205), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(G116), .B2(new_n205), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(G13), .A2(G33), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(G20), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n826), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n885), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n875), .B(new_n887), .C1(new_n776), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n822), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n825), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT102), .Z(G396));
  NOR2_X1   g0693(.A1(new_n506), .A2(new_n756), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n756), .A2(new_n416), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n424), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n896), .B2(new_n506), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(new_n816), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(new_n807), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n822), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n843), .A2(new_n263), .B1(new_n853), .B2(new_n215), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n289), .B1(new_n850), .B2(new_n213), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n838), .A2(G143), .B1(G150), .B2(new_n846), .ZN(new_n903));
  INV_X1    g0703(.A(G137), .ZN(new_n904));
  INV_X1    g0704(.A(new_n857), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .C1(new_n830), .C2(new_n836), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT34), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n901), .B(new_n902), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(G132), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n908), .B1(new_n907), .B2(new_n906), .C1(new_n909), .C2(new_n829), .ZN(new_n910));
  INV_X1    g0710(.A(new_n846), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n209), .A2(new_n836), .B1(new_n911), .B2(new_n863), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(new_n510), .C2(new_n905), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n865), .A2(G107), .B1(new_n854), .B2(G87), .ZN(new_n918));
  INV_X1    g0718(.A(G294), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n918), .B1(new_n860), .B2(new_n829), .C1(new_n839), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n287), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n910), .B1(new_n923), .B2(new_n844), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n826), .A2(new_n883), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n924), .A2(new_n826), .B1(new_n334), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n890), .C1(new_n884), .C2(new_n897), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n900), .A2(new_n927), .ZN(G384));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n459), .B1(new_n465), .B2(new_n215), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT16), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n318), .A3(new_n466), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(new_n457), .B1(new_n494), .B2(new_n752), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n443), .A2(new_n477), .A3(KEYINPUT85), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n487), .B1(new_n482), .B2(new_n486), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(KEYINPUT108), .A3(KEYINPUT37), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT108), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n934), .B1(new_n478), .B2(new_n488), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT37), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n494), .A2(new_n752), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n477), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n942), .B(new_n945), .C1(new_n936), .C2(new_n937), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n933), .A2(new_n457), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n501), .A2(new_n753), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(KEYINPUT38), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT38), .B1(new_n947), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n755), .A2(new_n351), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n390), .A2(new_n393), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n383), .B2(new_n389), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT107), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n712), .A2(new_n959), .A3(new_n954), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n707), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n962), .A2(new_n760), .A3(new_n772), .A4(new_n755), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n801), .A2(new_n756), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT31), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n801), .A2(KEYINPUT31), .A3(new_n756), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n897), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n929), .B1(new_n953), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n486), .A2(new_n752), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n501), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n498), .A2(new_n945), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n946), .B1(new_n942), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT38), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n950), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n897), .A2(new_n968), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT40), .A4(new_n961), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n970), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n331), .A2(new_n390), .A3(new_n424), .A4(new_n393), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n982), .A2(new_n501), .A3(new_n507), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n968), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n981), .B(new_n984), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(G330), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT39), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n947), .A2(new_n949), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n976), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(KEYINPUT39), .A3(new_n950), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n390), .A2(new_n756), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n897), .A2(new_n816), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n894), .B(KEYINPUT106), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n961), .C1(new_n951), .C2(new_n952), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n495), .A2(new_n496), .A3(new_n752), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n993), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(KEYINPUT29), .B(new_n756), .C1(new_n728), .C2(new_n740), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n983), .B1(new_n1000), .B2(new_n815), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n717), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n999), .B(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n986), .B(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n203), .B2(new_n748), .ZN(new_n1005));
  OAI21_X1  g0805(.A(G77), .B1(new_n263), .B2(new_n215), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1006), .A2(new_n223), .B1(G50), .B2(new_n215), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(G1), .A3(new_n747), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n209), .B1(new_n642), .B2(KEYINPUT35), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n222), .C1(KEYINPUT35), .C2(new_n642), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1005), .A2(new_n1008), .A3(new_n1012), .ZN(G367));
  NAND2_X1  g0813(.A1(new_n758), .A2(new_n759), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n760), .A2(new_n761), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n763), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n653), .B(new_n660), .C1(new_n646), .C2(new_n755), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n756), .A2(new_n734), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT42), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT42), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n765), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1018), .A2(new_n613), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1025), .A2(new_n660), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1024), .C1(new_n756), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n755), .B1(new_n686), .B2(new_n669), .ZN(new_n1028));
  MUX2_X1   g0828(.A(new_n720), .B(new_n719), .S(new_n1028), .Z(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT43), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n778), .A3(new_n1020), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1029), .A2(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n778), .A2(new_n1020), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1027), .A2(new_n1034), .A3(new_n1030), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n784), .B(KEYINPUT41), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n766), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n1020), .C1(new_n762), .C2(new_n764), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT45), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT44), .B1(new_n767), .B2(new_n1020), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT44), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n1021), .C1(new_n765), .C2(new_n766), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n779), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n778), .B1(new_n1049), .B2(new_n1043), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n823), .B1(new_n765), .B2(KEYINPUT109), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT109), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1017), .A2(new_n1052), .A3(new_n777), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1016), .B2(new_n763), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n762), .A4(new_n764), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1048), .A2(new_n1050), .A3(new_n1057), .A4(new_n819), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1040), .B1(new_n1058), .B2(new_n819), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n821), .A2(G1), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT110), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1038), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n911), .A2(new_n919), .B1(new_n853), .B2(new_n548), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT111), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n850), .B2(new_n209), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(KEYINPUT46), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT46), .B2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n287), .B1(new_n905), .B2(new_n860), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G303), .B2(new_n838), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n863), .B2(new_n836), .C1(new_n867), .C2(new_n829), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1067), .B(new_n1070), .C1(G107), .C2(new_n842), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n865), .A2(G58), .ZN(new_n1072));
  INV_X1    g0872(.A(G150), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n289), .B1(new_n904), .B2(new_n829), .C1(new_n839), .C2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n846), .A2(G159), .B1(new_n842), .B2(G68), .ZN(new_n1075));
  INV_X1    g0875(.A(G143), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n905), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n836), .A2(new_n213), .B1(new_n334), .B2(new_n853), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1071), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n822), .B1(new_n1082), .B2(new_n826), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n230), .A2(new_n876), .B1(new_n783), .B2(new_n408), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n886), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n888), .C2(new_n1029), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1062), .A2(new_n1086), .ZN(G387));
  NAND2_X1  g0887(.A1(new_n1057), .A2(new_n819), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1055), .A2(new_n818), .A3(new_n1056), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n784), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n838), .A2(G317), .B1(G311), .B2(new_n846), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n510), .B2(new_n836), .C1(new_n861), .C2(new_n905), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT48), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n863), .B2(new_n843), .C1(new_n919), .C2(new_n850), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n872), .A2(G326), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n289), .B1(new_n854), .B2(G116), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n289), .B1(new_n853), .B2(new_n544), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n842), .A2(new_n408), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n334), .B2(new_n850), .C1(new_n905), .C2(new_n830), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G50), .C2(new_n838), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n836), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1105), .A2(G68), .B1(new_n447), .B2(new_n846), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT114), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n1073), .C2(new_n829), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n237), .A2(new_n877), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT113), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(KEYINPUT113), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n781), .B1(G68), .B2(G77), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n406), .A2(G50), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT50), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n877), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1111), .A2(new_n876), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(G107), .B2(new_n205), .C1(new_n782), .C2(new_n881), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1109), .A2(new_n826), .B1(new_n886), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n762), .A2(new_n885), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1119), .A2(new_n890), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1090), .A2(new_n1122), .ZN(G393));
  OAI22_X1  g0923(.A1(new_n836), .A2(new_n406), .B1(new_n851), .B2(new_n853), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n911), .A2(new_n213), .B1(new_n215), .B2(new_n850), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n289), .B1(new_n829), .B2(new_n1076), .ZN(new_n1126));
  OR3_X1    g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT51), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n839), .A2(new_n830), .B1(new_n1073), .B2(new_n905), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n1128), .B2(new_n1129), .C1(new_n334), .C2(new_n843), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n838), .A2(G311), .B1(G317), .B2(new_n857), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT52), .Z(new_n1133));
  OAI22_X1  g0933(.A1(new_n836), .A2(new_n919), .B1(new_n585), .B2(new_n853), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n911), .A2(new_n510), .B1(new_n863), .B2(new_n850), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n287), .B1(new_n829), .B2(new_n861), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1133), .B(new_n1137), .C1(new_n209), .C2(new_n843), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n822), .B1(new_n1139), .B2(new_n826), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n876), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n886), .B1(new_n205), .B2(new_n548), .C1(new_n247), .C2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n888), .C2(new_n1020), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1061), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n785), .B1(new_n1144), .B2(new_n1088), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1058), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G390));
  NAND2_X1  g0949(.A1(new_n988), .A2(new_n991), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n992), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n995), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n816), .B2(new_n897), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n417), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT77), .B1(new_n405), .B2(new_n417), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n421), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n895), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1161), .A2(new_n506), .A3(new_n755), .A4(new_n814), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n995), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n961), .B1(new_n950), .B2(new_n977), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1151), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n963), .A2(new_n966), .A3(new_n806), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n506), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n894), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(G330), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT115), .B1(new_n1169), .B2(new_n1154), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT115), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n807), .A2(new_n1171), .A3(new_n897), .A4(new_n961), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1156), .A2(new_n1165), .A3(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1150), .A2(new_n1155), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n961), .A2(new_n897), .A3(G330), .A4(new_n968), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1175), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n425), .A2(G330), .A3(new_n968), .A4(new_n508), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n717), .B(new_n1180), .C1(new_n817), .C2(new_n509), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT116), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT116), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1001), .A2(new_n1183), .A3(new_n717), .A4(new_n1180), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n897), .A2(G330), .A3(new_n968), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1163), .B1(new_n1154), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1169), .A2(new_n1154), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1177), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n996), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT117), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1173), .A2(new_n1187), .B1(new_n1190), .B2(new_n996), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT117), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1179), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1185), .A2(new_n1192), .A3(KEYINPUT117), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1196), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1156), .A2(new_n1165), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1177), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .A4(new_n1175), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n784), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT118), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1198), .A2(new_n1203), .A3(new_n1206), .A4(new_n784), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1179), .A2(new_n1061), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1150), .A2(new_n883), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n850), .A2(new_n1073), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT53), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n213), .B2(new_n853), .C1(new_n904), .C2(new_n911), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n289), .B1(new_n830), .B2(new_n843), .C1(new_n839), .C2(new_n909), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT54), .B(G143), .Z(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1105), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(new_n829), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1213), .B(new_n1218), .C1(G128), .C2(new_n857), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n289), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT119), .B1(new_n852), .B2(new_n289), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n857), .A2(G283), .B1(new_n842), .B2(G77), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n838), .A2(G116), .B1(G68), .B2(new_n854), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n919), .B2(new_n829), .C1(new_n548), .C2(new_n836), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G107), .C2(new_n846), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n826), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n444), .A2(new_n925), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1210), .A2(new_n890), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1209), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1208), .A2(new_n1230), .ZN(G378));
  INV_X1    g1031(.A(KEYINPUT55), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n331), .B(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n327), .A2(new_n752), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT56), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1233), .B(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n883), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n850), .A2(new_n334), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n853), .A2(new_n263), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G116), .C2(new_n857), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n215), .B2(new_n843), .C1(new_n544), .C2(new_n911), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G41), .B1(new_n872), .B2(G283), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n409), .B2(new_n836), .C1(new_n839), .C2(new_n585), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1241), .A2(new_n289), .A3(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT120), .Z(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n865), .A2(new_n1215), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n843), .B2(new_n1073), .C1(new_n905), .C2(new_n1217), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n838), .A2(G128), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n904), .B2(new_n836), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(G132), .C2(new_n846), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT59), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G41), .B1(new_n854), .B2(G159), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G33), .B1(new_n872), .B2(G124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n280), .A2(new_n278), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n213), .B1(new_n1257), .B2(G41), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1246), .A2(new_n1247), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1259), .A2(new_n826), .B1(new_n213), .B2(new_n925), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1237), .A2(new_n890), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n969), .B1(new_n990), .B2(new_n950), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G330), .B(new_n980), .C1(new_n1263), .C2(KEYINPUT40), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1236), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1236), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n970), .A2(G330), .A3(new_n1266), .A4(new_n980), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n999), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n999), .A3(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1262), .B1(new_n1272), .B2(new_n1061), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1198), .A2(new_n1185), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1274), .B2(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1195), .B1(new_n1276), .B2(new_n1179), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1265), .A2(new_n999), .A3(new_n1267), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n999), .B1(new_n1267), .B2(new_n1265), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT57), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n784), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1273), .B1(new_n1275), .B2(new_n1281), .ZN(G375));
  OAI221_X1 g1082(.A(new_n1102), .B1(new_n544), .B2(new_n850), .C1(new_n905), .C2(new_n919), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n287), .B1(new_n334), .B2(new_n853), .C1(new_n839), .C2(new_n863), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1105), .A2(G107), .B1(G116), .B2(new_n846), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1283), .B(new_n1284), .C1(KEYINPUT122), .C2(new_n1285), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1286), .B1(KEYINPUT122), .B2(new_n1285), .C1(new_n510), .C2(new_n829), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n843), .A2(new_n213), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n905), .A2(new_n909), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1289), .A2(KEYINPUT123), .B1(new_n836), .B2(new_n1073), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(KEYINPUT123), .B2(new_n1289), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n846), .A2(new_n1215), .B1(new_n865), .B2(G159), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n287), .B1(new_n872), .B2(G128), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1239), .B1(new_n838), .B2(G137), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1287), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1296), .A2(new_n826), .B1(new_n215), .B2(new_n925), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n890), .C1(new_n961), .C2(new_n884), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1194), .B2(new_n1145), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT121), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT121), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1200), .A3(new_n1199), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1300), .B1(new_n1306), .B2(new_n1040), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1307), .A2(KEYINPUT124), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(KEYINPUT124), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(G381));
  INV_X1    g1110(.A(G381), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1204), .A2(new_n1230), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(G375), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1062), .A2(new_n1086), .A3(new_n1148), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1311), .A2(new_n1312), .A3(new_n1314), .A4(new_n1316), .ZN(G407));
  INV_X1    g1117(.A(new_n1314), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G407), .B(G213), .C1(G343), .C2(new_n1318), .ZN(G409));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  INV_X1    g1121(.A(G384), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT60), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT60), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n785), .B(new_n1324), .C1(new_n1325), .C2(new_n1305), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1322), .B1(new_n1326), .B2(new_n1299), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT60), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1304), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT121), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n784), .B(new_n1323), .C1(new_n1328), .C2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(G384), .A3(new_n1300), .ZN(new_n1333));
  INV_X1    g1133(.A(G213), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(G343), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(G2897), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1327), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1336), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1324), .B1(new_n1325), .B2(new_n1305), .ZN(new_n1339));
  AOI211_X1 g1139(.A(new_n1322), .B(new_n1299), .C1(new_n1339), .C2(new_n784), .ZN(new_n1340));
  AOI21_X1  g1140(.A(G384), .B1(new_n1332), .B2(new_n1300), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1338), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  AOI22_X1  g1142(.A1(new_n1200), .A2(new_n1199), .B1(new_n1202), .B2(new_n1175), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1272), .B(new_n1039), .C1(new_n1343), .C2(new_n1195), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1313), .B1(new_n1273), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1273), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT57), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1347), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n785), .B1(new_n1274), .B2(new_n1348), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1277), .B2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1346), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1345), .B1(G378), .B2(new_n1352), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1337), .B(new_n1342), .C1(new_n1353), .C2(new_n1335), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1344), .A2(new_n1273), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1355), .A2(new_n1230), .A3(new_n1204), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1230), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1357), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1356), .B1(G375), .B2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1335), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1321), .B1(new_n1354), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1321), .ZN(new_n1364));
  AND2_X1   g1164(.A1(G393), .A2(G396), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(G393), .A2(G396), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G387), .A2(G390), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1368), .B2(new_n1315), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1368), .A2(new_n1315), .A3(new_n1367), .ZN(new_n1371));
  AOI21_X1  g1171(.A(KEYINPUT61), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1364), .A2(new_n1372), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1320), .B1(new_n1363), .B2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1342), .A2(new_n1337), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1375), .B1(new_n1361), .B2(new_n1359), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1359), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1377));
  OAI21_X1  g1177(.A(KEYINPUT63), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT61), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1367), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1148), .B1(new_n1062), .B2(new_n1086), .ZN(new_n1381));
  NOR3_X1   g1181(.A1(new_n1316), .A2(new_n1380), .A3(new_n1381), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1379), .B1(new_n1382), .B2(new_n1369), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1383), .B1(new_n1321), .B2(new_n1362), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1378), .A2(KEYINPUT125), .A3(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1374), .A2(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT62), .ZN(new_n1387));
  OAI21_X1  g1187(.A(new_n1387), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1362), .A2(KEYINPUT62), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1388), .A2(new_n1379), .A3(new_n1389), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1382), .A2(new_n1369), .ZN(new_n1391));
  XOR2_X1   g1191(.A(new_n1391), .B(KEYINPUT126), .Z(new_n1392));
  NAND2_X1  g1192(.A1(new_n1390), .A2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1386), .A2(new_n1393), .ZN(G405));
  XNOR2_X1  g1194(.A(new_n1360), .B(KEYINPUT127), .ZN(new_n1395));
  NOR2_X1   g1195(.A1(new_n1352), .A2(new_n1313), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1396), .B1(G378), .B2(new_n1352), .ZN(new_n1397));
  XNOR2_X1  g1197(.A(new_n1395), .B(new_n1397), .ZN(new_n1398));
  INV_X1    g1198(.A(new_n1391), .ZN(new_n1399));
  XNOR2_X1  g1199(.A(new_n1398), .B(new_n1399), .ZN(G402));
endmodule


