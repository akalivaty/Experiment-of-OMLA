

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n727), .ZN(n690) );
  NAND2_X2 U553 ( .A1(n679), .A2(n764), .ZN(n727) );
  XNOR2_X1 U554 ( .A(n525), .B(KEYINPUT92), .ZN(G164) );
  NOR2_X1 U555 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  INV_X1 U557 ( .A(KEYINPUT31), .ZN(n722) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n758), .ZN(n739) );
  AND2_X1 U559 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U560 ( .A1(n799), .A2(n798), .ZN(n801) );
  NOR2_X1 U561 ( .A1(n628), .A2(G651), .ZN(n647) );
  AND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n869) );
  NAND2_X1 U563 ( .A1(G114), .A2(n869), .ZN(n517) );
  INV_X1 U564 ( .A(G2105), .ZN(n519) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n519), .ZN(n870) );
  NAND2_X1 U566 ( .A1(G126), .A2(n870), .ZN(n516) );
  NAND2_X1 U567 ( .A1(n517), .A2(n516), .ZN(n524) );
  XOR2_X1 U568 ( .A(KEYINPUT17), .B(n518), .Z(n873) );
  NAND2_X1 U569 ( .A1(n873), .A2(G138), .ZN(n522) );
  AND2_X1 U570 ( .A1(G2104), .A2(n519), .ZN(n520) );
  XNOR2_X2 U571 ( .A(n520), .B(KEYINPUT64), .ZN(n875) );
  NAND2_X1 U572 ( .A1(G102), .A2(n875), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U575 ( .A1(G101), .A2(n875), .ZN(n526) );
  XOR2_X1 U576 ( .A(n526), .B(KEYINPUT23), .Z(n528) );
  NAND2_X1 U577 ( .A1(n870), .A2(G125), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT65), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G137), .A2(n873), .ZN(n530) );
  AND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n869), .A2(G113), .ZN(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT66), .B(n532), .ZN(n533) );
  AND2_X2 U584 ( .A1(n534), .A2(n533), .ZN(G160) );
  XNOR2_X1 U585 ( .A(KEYINPUT9), .B(KEYINPUT73), .ZN(n539) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n628) );
  XNOR2_X1 U587 ( .A(KEYINPUT67), .B(G651), .ZN(n541) );
  NOR2_X1 U588 ( .A1(n628), .A2(n541), .ZN(n535) );
  XNOR2_X1 U589 ( .A(KEYINPUT68), .B(n535), .ZN(n640) );
  NAND2_X1 U590 ( .A1(G77), .A2(n640), .ZN(n537) );
  NOR2_X1 U591 ( .A1(G543), .A2(G651), .ZN(n641) );
  NAND2_X1 U592 ( .A1(G90), .A2(n641), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n539), .B(n538), .ZN(n546) );
  NAND2_X1 U595 ( .A1(n647), .A2(G52), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT72), .ZN(n544) );
  NOR2_X1 U597 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n542), .Z(n645) );
  NAND2_X1 U599 ( .A1(G64), .A2(n645), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n546), .A2(n545), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  NAND2_X1 U604 ( .A1(n647), .A2(G51), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G63), .A2(n645), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n549), .Z(n557) );
  NAND2_X1 U608 ( .A1(n640), .A2(G76), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT81), .B(n550), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n641), .A2(G89), .ZN(n551) );
  XOR2_X1 U611 ( .A(n551), .B(KEYINPUT4), .Z(n552) );
  NOR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U613 ( .A(KEYINPUT5), .B(n554), .Z(n555) );
  XNOR2_X1 U614 ( .A(KEYINPUT82), .B(n555), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U616 ( .A(KEYINPUT7), .B(n558), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n819) );
  NAND2_X1 U621 ( .A1(n819), .A2(G567), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n560), .B(KEYINPUT77), .ZN(n561) );
  XNOR2_X1 U623 ( .A(KEYINPUT11), .B(n561), .ZN(G234) );
  XOR2_X1 U624 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n563) );
  NAND2_X1 U625 ( .A1(G56), .A2(n645), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n570) );
  XNOR2_X1 U627 ( .A(KEYINPUT79), .B(KEYINPUT13), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n641), .A2(G81), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G68), .A2(n640), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n647), .A2(G43), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n967) );
  INV_X1 U636 ( .A(G860), .ZN(n592) );
  OR2_X1 U637 ( .A1(n967), .A2(n592), .ZN(G153) );
  XOR2_X1 U638 ( .A(G171), .B(KEYINPUT80), .Z(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n641), .A2(G92), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G66), .A2(n645), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G79), .A2(n640), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G54), .A2(n647), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT15), .B(n579), .Z(n964) );
  OR2_X1 U648 ( .A1(n964), .A2(G868), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G78), .A2(n640), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G91), .A2(n641), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT74), .B(n584), .Z(n588) );
  NAND2_X1 U654 ( .A1(n645), .A2(G65), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n647), .A2(G53), .ZN(n585) );
  AND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(G299) );
  XNOR2_X1 U658 ( .A(KEYINPUT83), .B(G868), .ZN(n589) );
  NOR2_X1 U659 ( .A1(G286), .A2(n589), .ZN(n591) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n593), .A2(n964), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n967), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G868), .A2(n964), .ZN(n595) );
  NOR2_X1 U667 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT84), .B(n598), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G111), .A2(n869), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G99), .A2(n875), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT85), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G135), .A2(n873), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n870), .A2(G123), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n990) );
  XNOR2_X1 U679 ( .A(n990), .B(G2096), .ZN(n608) );
  INV_X1 U680 ( .A(G2100), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G156) );
  NAND2_X1 U682 ( .A1(n964), .A2(G559), .ZN(n659) );
  XNOR2_X1 U683 ( .A(n967), .B(n659), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n609), .A2(G860), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G80), .A2(n640), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G93), .A2(n641), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U688 ( .A(KEYINPUT86), .B(n612), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n647), .A2(G55), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G67), .A2(n645), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n662) );
  XOR2_X1 U693 ( .A(n617), .B(n662), .Z(G145) );
  NAND2_X1 U694 ( .A1(G86), .A2(n641), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G48), .A2(n647), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n640), .A2(G73), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT2), .B(n620), .Z(n621) );
  NOR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G61), .A2(n645), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(G305) );
  NAND2_X1 U702 ( .A1(G49), .A2(n647), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n645), .A2(n627), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G87), .A2(n628), .ZN(n629) );
  XOR2_X1 U707 ( .A(KEYINPUT87), .B(n629), .Z(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G75), .A2(n640), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G88), .A2(n641), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U712 ( .A(KEYINPUT89), .B(n634), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n647), .A2(G50), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G62), .A2(n645), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT88), .B(n637), .Z(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(G303) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G72), .A2(n640), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G85), .A2(n641), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(n644), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n645), .A2(G60), .ZN(n646) );
  XOR2_X1 U724 ( .A(KEYINPUT70), .B(n646), .Z(n650) );
  NAND2_X1 U725 ( .A1(G47), .A2(n647), .ZN(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT71), .B(n648), .ZN(n649) );
  NOR2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(G290) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(G305), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(n662), .ZN(n656) );
  INV_X1 U732 ( .A(G299), .ZN(n689) );
  XNOR2_X1 U733 ( .A(n689), .B(G166), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(n967), .ZN(n893) );
  XOR2_X1 U737 ( .A(n893), .B(n659), .Z(n660) );
  NAND2_X1 U738 ( .A1(G868), .A2(n660), .ZN(n664) );
  INV_X1 U739 ( .A(G868), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT76), .B(G82), .Z(G220) );
  XNOR2_X1 U749 ( .A(KEYINPUT75), .B(G132), .ZN(G219) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U752 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n671), .A2(G96), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n672), .A2(G218), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(KEYINPUT91), .ZN(n825) );
  NAND2_X1 U756 ( .A1(n825), .A2(G2106), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U758 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G108), .A2(n675), .ZN(n826) );
  NAND2_X1 U760 ( .A1(n826), .A2(G567), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n827) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n827), .A2(n678), .ZN(n824) );
  NAND2_X1 U764 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n763) );
  INV_X1 U766 ( .A(n763), .ZN(n679) );
  NOR2_X1 U767 ( .A1(G1384), .A2(G164), .ZN(n764) );
  NAND2_X2 U768 ( .A1(G8), .A2(n727), .ZN(n758) );
  NOR2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n745) );
  NAND2_X1 U770 ( .A1(n745), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U771 ( .A1(n758), .A2(n680), .ZN(n750) );
  OR2_X1 U772 ( .A1(n690), .A2(G1961), .ZN(n682) );
  XNOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .ZN(n939) );
  NAND2_X1 U774 ( .A1(n690), .A2(n939), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n719) );
  NAND2_X1 U776 ( .A1(G171), .A2(n719), .ZN(n683) );
  XNOR2_X1 U777 ( .A(KEYINPUT100), .B(n683), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n690), .A2(G2072), .ZN(n684) );
  XNOR2_X1 U779 ( .A(n684), .B(KEYINPUT27), .ZN(n686) );
  INV_X1 U780 ( .A(G1956), .ZN(n914) );
  NOR2_X1 U781 ( .A1(n914), .A2(n690), .ZN(n685) );
  NOR2_X1 U782 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n687) );
  XOR2_X1 U784 ( .A(n687), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n707) );
  NOR2_X1 U786 ( .A1(n690), .A2(G1348), .ZN(n692) );
  NOR2_X1 U787 ( .A1(G2067), .A2(n727), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n699) );
  INV_X1 U789 ( .A(G1996), .ZN(n940) );
  NOR2_X1 U790 ( .A1(n763), .A2(n940), .ZN(n693) );
  AND2_X1 U791 ( .A1(n764), .A2(n693), .ZN(n694) );
  XOR2_X1 U792 ( .A(n694), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U793 ( .A1(n727), .A2(G1341), .ZN(n695) );
  AND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U795 ( .A(n967), .ZN(n702) );
  AND2_X1 U796 ( .A1(n702), .A2(n964), .ZN(n697) );
  NAND2_X1 U797 ( .A1(n701), .A2(n697), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U799 ( .A(KEYINPUT101), .B(n700), .Z(n705) );
  AND2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U801 ( .A1(n964), .A2(n703), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n711) );
  XOR2_X1 U805 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n710) );
  XNOR2_X1 U806 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n725) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n727), .ZN(n736) );
  NOR2_X1 U809 ( .A1(n739), .A2(n736), .ZN(n715) );
  INV_X1 U810 ( .A(KEYINPUT103), .ZN(n714) );
  XNOR2_X1 U811 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n716), .A2(G8), .ZN(n717) );
  XNOR2_X1 U813 ( .A(n717), .B(KEYINPUT30), .ZN(n718) );
  NOR2_X1 U814 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U815 ( .A1(G171), .A2(n719), .ZN(n720) );
  XNOR2_X1 U816 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n737) );
  NAND2_X1 U818 ( .A1(n737), .A2(G286), .ZN(n734) );
  INV_X1 U819 ( .A(G8), .ZN(n732) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n758), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n726), .B(KEYINPUT104), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n727), .A2(G2090), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n735), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U827 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U828 ( .A(n737), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n754) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n971) );
  NAND2_X1 U834 ( .A1(n754), .A2(n971), .ZN(n746) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NAND2_X1 U836 ( .A1(n746), .A2(n965), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n747), .A2(n758), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n976) );
  NAND2_X1 U841 ( .A1(n751), .A2(n976), .ZN(n762) );
  NOR2_X1 U842 ( .A1(G2090), .A2(G303), .ZN(n752) );
  NAND2_X1 U843 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U845 ( .A1(n755), .A2(n758), .ZN(n760) );
  NOR2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XOR2_X1 U847 ( .A(n756), .B(KEYINPUT24), .Z(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n799) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n814) );
  NAND2_X1 U852 ( .A1(n873), .A2(G140), .ZN(n765) );
  XOR2_X1 U853 ( .A(KEYINPUT93), .B(n765), .Z(n767) );
  NAND2_X1 U854 ( .A1(G104), .A2(n875), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U856 ( .A(KEYINPUT34), .B(n768), .ZN(n775) );
  NAND2_X1 U857 ( .A1(n870), .A2(G128), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT94), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G116), .A2(n869), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(KEYINPUT95), .B(n772), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT35), .B(n773), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT36), .ZN(n777) );
  XOR2_X1 U865 ( .A(n777), .B(KEYINPUT96), .Z(n857) );
  XOR2_X1 U866 ( .A(KEYINPUT37), .B(G2067), .Z(n811) );
  AND2_X1 U867 ( .A1(n857), .A2(n811), .ZN(n1002) );
  NAND2_X1 U868 ( .A1(n814), .A2(n1002), .ZN(n808) );
  NAND2_X1 U869 ( .A1(G117), .A2(n869), .ZN(n779) );
  NAND2_X1 U870 ( .A1(G129), .A2(n870), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n875), .A2(G105), .ZN(n780) );
  XOR2_X1 U873 ( .A(KEYINPUT97), .B(n780), .Z(n781) );
  XNOR2_X1 U874 ( .A(n781), .B(KEYINPUT38), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G141), .A2(n873), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U878 ( .A(KEYINPUT98), .B(n786), .Z(n856) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n856), .ZN(n787) );
  XNOR2_X1 U880 ( .A(n787), .B(KEYINPUT99), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n873), .A2(G131), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G95), .A2(n875), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G107), .A2(n869), .ZN(n791) );
  NAND2_X1 U885 ( .A1(G119), .A2(n870), .ZN(n790) );
  NAND2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n885) );
  AND2_X1 U888 ( .A1(G1991), .A2(n885), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n1000) );
  INV_X1 U890 ( .A(n814), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n1000), .A2(n796), .ZN(n804) );
  INV_X1 U892 ( .A(n804), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n808), .A2(n797), .ZN(n798) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U895 ( .A1(n982), .A2(n814), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n817) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n856), .ZN(n995) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n885), .ZN(n991) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U900 ( .A1(n991), .A2(n802), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT105), .B(n805), .Z(n806) );
  NOR2_X1 U903 ( .A1(n995), .A2(n806), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT106), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n857), .A2(n811), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT107), .ZN(n1004) );
  NAND2_X1 U909 ( .A1(n813), .A2(n1004), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n819), .ZN(G217) );
  NAND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n821) );
  INV_X1 U915 ( .A(G661), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n827), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2474), .B(G1976), .Z(n829) );
  XNOR2_X1 U928 ( .A(G1956), .B(G1961), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U930 ( .A(n830), .B(KEYINPUT112), .Z(n832) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(G1981), .B(G1971), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1966), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2678), .Z(n840) );
  XNOR2_X1 U940 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2096), .B(G2100), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U948 ( .A(G2078), .B(G2084), .Z(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G227) );
  NAND2_X1 U950 ( .A1(G124), .A2(n870), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n869), .A2(G112), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n873), .A2(G136), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G100), .A2(n875), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U957 ( .A1(n855), .A2(n854), .ZN(G162) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n868) );
  NAND2_X1 U959 ( .A1(n873), .A2(G139), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G103), .A2(n875), .ZN(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n870), .A2(G127), .ZN(n860) );
  XNOR2_X1 U963 ( .A(KEYINPUT115), .B(n860), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n869), .A2(G115), .ZN(n861) );
  XOR2_X1 U965 ( .A(n861), .B(KEYINPUT116), .Z(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n864), .Z(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT117), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n1007) );
  XNOR2_X1 U970 ( .A(n868), .B(n1007), .ZN(n891) );
  NAND2_X1 U971 ( .A1(G118), .A2(n869), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G130), .A2(n870), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n873), .A2(G142), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT114), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G106), .A2(n875), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U980 ( .A(G160), .B(n881), .ZN(n889) );
  XOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n883) );
  XNOR2_X1 U982 ( .A(G162), .B(KEYINPUT118), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n990), .B(n884), .ZN(n887) );
  XOR2_X1 U985 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U989 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U990 ( .A(KEYINPUT119), .B(n893), .Z(n895) );
  XNOR2_X1 U991 ( .A(n964), .B(G286), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(G171), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2438), .B(KEYINPUT108), .Z(n899) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2430), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n900), .B(G2435), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2446), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G20), .B(n914), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G1341), .B(G19), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(G1981), .B(G6), .ZN(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT59), .B(G1348), .Z(n919) );
  XNOR2_X1 U1021 ( .A(G4), .B(n919), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT60), .B(n922), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT126), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G21), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(G1961), .B(G5), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G23), .B(G1976), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1032 ( .A(G1986), .B(G24), .Z(n930) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n932), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT61), .B(n935), .Z(n936) );
  NOR2_X1 U1037 ( .A1(G16), .A2(n936), .ZN(n963) );
  XOR2_X1 U1038 ( .A(G2090), .B(G35), .Z(n953) );
  XOR2_X1 U1039 ( .A(G1991), .B(G25), .Z(n937) );
  NAND2_X1 U1040 ( .A1(n937), .A2(G28), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(KEYINPUT122), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G27), .B(n939), .ZN(n946) );
  XOR2_X1 U1043 ( .A(G2067), .B(G26), .Z(n942) );
  XNOR2_X1 U1044 ( .A(n940), .B(G32), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(n950), .B(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT53), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(G34), .B(G2084), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(KEYINPUT55), .B(n957), .ZN(n959) );
  INV_X1 U1058 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(G11), .ZN(n961) );
  XOR2_X1 U1061 ( .A(KEYINPUT125), .B(n961), .Z(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n988) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1064 ( .A(n964), .B(G1348), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1070 ( .A(G171), .B(G1961), .Z(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n978), .Z(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G1956), .B(G299), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT127), .ZN(n1018) );
  XNOR2_X1 U1083 ( .A(G160), .B(G2084), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n998) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT51), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT120), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G2078), .B(KEYINPUT121), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(G164), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1007), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1010), .Z(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

