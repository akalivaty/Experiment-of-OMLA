//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n192), .A2(KEYINPUT64), .A3(G146), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT64), .B1(new_n192), .B2(G146), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n189), .B(new_n191), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(G143), .B2(new_n188), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n199), .B2(new_n190), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI211_X1 g025(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n202), .C2(G134), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n206), .B(new_n207), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT67), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT68), .B(new_n201), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n189), .B(new_n220), .C1(new_n193), .C2(new_n194), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n197), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n226), .B2(new_n213), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  AOI211_X1 g043(.A(new_n229), .B(new_n224), .C1(new_n226), .C2(new_n213), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n218), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n213), .A2(new_n215), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(new_n236), .B2(new_n201), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n239), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n224), .ZN(new_n250));
  INV_X1    g064(.A(new_n213), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n210), .B1(new_n204), .B2(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n209), .A2(new_n208), .A3(new_n210), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n207), .B1(new_n255), .B2(new_n206), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n250), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n201), .A2(new_n213), .A3(new_n215), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(KEYINPUT30), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT69), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n238), .A2(new_n249), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT26), .B(G101), .Z(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n262), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n201), .A2(new_n213), .A3(new_n215), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n227), .A2(new_n270), .A3(new_n249), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n249), .B1(new_n231), .B2(new_n237), .ZN(new_n276));
  INV_X1    g090(.A(new_n249), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n257), .A2(new_n277), .A3(new_n258), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n278), .A2(KEYINPUT71), .A3(new_n275), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT71), .B1(new_n278), .B2(new_n275), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n269), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n261), .A2(new_n285), .A3(new_n272), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n274), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n280), .B2(new_n281), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n271), .B2(KEYINPUT28), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n278), .A2(KEYINPUT71), .A3(new_n275), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n277), .B1(new_n257), .B2(new_n258), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n271), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT29), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n201), .B1(new_n216), .B2(new_n217), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n257), .A2(new_n229), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n309), .A3(new_n218), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n271), .B1(new_n310), .B2(new_n249), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n303), .B(new_n282), .C1(new_n311), .C2(new_n275), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n302), .A2(new_n268), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n261), .A2(new_n303), .A3(new_n278), .A4(new_n269), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G472), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n291), .A2(new_n292), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n263), .A2(new_n264), .A3(G214), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n192), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n263), .A2(new_n264), .A3(G143), .A4(G214), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT17), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(KEYINPUT90), .A3(G131), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n207), .A3(new_n321), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G125), .A3(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n331), .B2(G140), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n335), .A2(new_n188), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n188), .B1(new_n335), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n325), .A2(new_n327), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n329), .B(new_n340), .C1(new_n341), .C2(new_n326), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT18), .A2(G131), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n322), .B(new_n346), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n333), .A2(G125), .A3(G140), .ZN(new_n348));
  AOI21_X1  g162(.A(G140), .B1(new_n333), .B2(G125), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT89), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n351), .A3(new_n334), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(G146), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n188), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n342), .A2(new_n345), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n341), .A2(new_n328), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT19), .A4(new_n352), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n332), .A2(new_n351), .A3(new_n334), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n351), .B1(new_n332), .B2(new_n334), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT19), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n354), .B2(new_n364), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n361), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n339), .B1(new_n368), .B2(new_n188), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n350), .A2(KEYINPUT19), .A3(new_n352), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n366), .ZN(new_n373));
  AOI21_X1  g187(.A(G146), .B1(new_n373), .B2(new_n361), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(KEYINPUT92), .A3(new_n339), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n357), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n345), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n358), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G475), .A2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT93), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n188), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n335), .A2(new_n337), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G146), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n370), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT92), .B1(new_n374), .B2(new_n339), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n359), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n345), .B1(new_n388), .B2(new_n357), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n379), .B1(new_n389), .B2(new_n358), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT20), .ZN(new_n392));
  INV_X1    g206(.A(new_n390), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n382), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n345), .B1(new_n342), .B2(new_n357), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n315), .B1(new_n358), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G475), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT95), .B1(new_n190), .B2(G143), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT95), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n192), .A3(G128), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n192), .A2(G128), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(G134), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(G116), .B(G122), .Z(new_n406));
  OR2_X1    g220(.A1(KEYINPUT81), .A2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT81), .A2(G107), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n406), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n405), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n404), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n400), .A2(new_n402), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n413), .ZN(new_n418));
  OAI21_X1  g232(.A(G134), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n412), .B(new_n419), .C1(new_n411), .C2(new_n410), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n243), .A2(G122), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n406), .B2(KEYINPUT14), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n204), .B1(new_n417), .B2(new_n416), .ZN(new_n425));
  OAI221_X1 g239(.A(new_n424), .B1(new_n406), .B2(new_n409), .C1(new_n405), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n420), .A2(new_n426), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n315), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT97), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n315), .B(new_n264), .C1(G234), .C2(G237), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G952), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  INV_X1    g258(.A(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n263), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n438), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n396), .A2(new_n399), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT25), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n190), .A2(G119), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n241), .A2(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT24), .B(G110), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT73), .B1(new_n190), .B2(G119), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT73), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n459), .C1(new_n241), .C2(G128), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G110), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n457), .B(new_n464), .C1(new_n338), .C2(new_n339), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n241), .B2(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT23), .ZN(new_n467));
  INV_X1    g281(.A(G110), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n454), .A4(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n455), .A2(new_n456), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n355), .A3(new_n385), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT76), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n472), .A3(KEYINPUT76), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT75), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT22), .B(G137), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n465), .A2(new_n472), .A3(KEYINPUT76), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT76), .B1(new_n465), .B2(new_n472), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n451), .B(new_n452), .C1(new_n486), .C2(KEYINPUT77), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n429), .B1(G234), .B2(new_n315), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n483), .A2(new_n484), .A3(new_n480), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n473), .A2(new_n481), .A3(new_n474), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n315), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT78), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT25), .B1(new_n486), .B2(new_n451), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n487), .B(new_n488), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n452), .B1(new_n491), .B2(KEYINPUT78), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n451), .B1(new_n486), .B2(KEYINPUT77), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n500), .A2(KEYINPUT79), .A3(new_n487), .A4(new_n488), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n489), .A2(new_n490), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT80), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n488), .A2(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G469), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n199), .A2(new_n190), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n192), .A2(G146), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT64), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n188), .B2(G143), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n192), .A2(KEYINPUT64), .A3(G146), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n195), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n407), .A2(new_n516), .A3(G104), .A4(new_n408), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n421), .B1(new_n516), .B2(G104), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(G104), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G101), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(G104), .B2(G107), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n409), .B2(G104), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT10), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n517), .A2(new_n520), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(G101), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n521), .B1(new_n517), .B2(new_n520), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n250), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n251), .A2(new_n256), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n522), .A2(new_n524), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n201), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n527), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  INV_X1    g352(.A(G227), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n522), .A2(new_n524), .ZN(new_n544));
  OAI21_X1  g358(.A(G128), .B1(new_n510), .B2(new_n198), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n514), .A2(new_n191), .B1(new_n545), .B2(new_n197), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n525), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g363(.A(new_n534), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT84), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n525), .A2(new_n551), .A3(new_n547), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n226), .B2(new_n213), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT83), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n548), .A2(KEYINPUT83), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n543), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n527), .A2(new_n533), .A3(new_n536), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n550), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n542), .B1(new_n565), .B2(new_n537), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n508), .B(new_n315), .C1(new_n563), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n564), .A2(new_n550), .ZN(new_n569));
  INV_X1    g383(.A(new_n537), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n541), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n553), .A2(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n543), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT85), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n508), .A4(new_n315), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n525), .A2(new_n551), .A3(new_n547), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n551), .B1(new_n525), .B2(new_n547), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(new_n577), .A3(new_n534), .ZN(new_n578));
  INV_X1    g392(.A(new_n561), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT83), .B1(new_n548), .B2(new_n557), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n578), .A2(KEYINPUT12), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n542), .B1(new_n581), .B2(new_n537), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n569), .A2(new_n543), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n315), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n568), .A2(new_n575), .B1(new_n584), .B2(G469), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G214), .B1(G237), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n249), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n593));
  OAI21_X1  g407(.A(G113), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n593), .A2(new_n595), .B1(new_n245), .B2(new_n240), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n535), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(G110), .B(G122), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n592), .A2(new_n597), .A3(new_n599), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT86), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT6), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n195), .A2(new_n200), .A3(new_n331), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n331), .B1(new_n221), .B2(new_n223), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT87), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(KEYINPUT87), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G224), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n610), .B(new_n612), .C1(new_n613), .C2(G953), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(G953), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT87), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n224), .A2(G125), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n607), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n615), .B1(new_n618), .B2(new_n611), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n598), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n606), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT7), .ZN(new_n623));
  OAI22_X1  g437(.A1(new_n618), .A2(new_n611), .B1(new_n623), .B2(new_n615), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n599), .B(KEYINPUT8), .Z(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n596), .B2(new_n544), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n595), .A2(KEYINPUT88), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n594), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n593), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(new_n246), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n631), .B2(new_n544), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n615), .A2(new_n623), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n610), .A2(new_n612), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n624), .A2(new_n632), .A3(new_n634), .A4(new_n602), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n315), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n591), .B1(new_n622), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n606), .A2(new_n620), .A3(new_n621), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n315), .A3(new_n590), .A4(new_n635), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n589), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n585), .A2(new_n587), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n318), .A2(new_n450), .A3(new_n507), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  NAND2_X1  g458(.A1(new_n640), .A2(new_n447), .ZN(new_n645));
  INV_X1    g459(.A(new_n399), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT20), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n391), .B1(new_n390), .B2(KEYINPUT20), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n649), .B2(new_n395), .ZN(new_n650));
  NOR2_X1   g464(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n432), .B(new_n433), .C1(new_n651), .C2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n436), .A2(G902), .ZN(new_n655));
  INV_X1    g469(.A(new_n434), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n435), .A2(new_n436), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT99), .B1(new_n650), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n396), .B2(new_n399), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n645), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n287), .A2(new_n315), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n666), .A2(G472), .B1(new_n288), .B2(new_n287), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n568), .A2(new_n575), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n584), .A2(G469), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n587), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n667), .A2(new_n507), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  NAND2_X1  g488(.A1(new_n438), .A2(new_n399), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT100), .B1(new_n647), .B2(new_n648), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n382), .A2(new_n677), .A3(new_n392), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n395), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(new_n682), .A3(new_n395), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n675), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n447), .B(KEYINPUT102), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n640), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n671), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NOR2_X1   g503(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n473), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n504), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n497), .A2(new_n501), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n670), .A2(new_n640), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n450), .A3(new_n667), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT37), .B(G110), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT103), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n695), .B(new_n697), .ZN(G12));
  NAND2_X1  g512(.A1(new_n681), .A2(new_n683), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT32), .B1(new_n287), .B2(new_n288), .ZN(new_n701));
  INV_X1    g515(.A(G472), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n314), .A2(new_n315), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n302), .A2(new_n312), .A3(new_n268), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n700), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n670), .A2(new_n693), .A3(new_n640), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n675), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n446), .B(KEYINPUT104), .ZN(new_n710));
  INV_X1    g524(.A(G900), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n441), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n699), .A2(new_n708), .A3(new_n709), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G128), .ZN(G30));
  XOR2_X1   g530(.A(new_n713), .B(KEYINPUT39), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n670), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT40), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n718), .B(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n396), .A2(new_n399), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n637), .A2(new_n639), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT38), .Z(new_n727));
  INV_X1    g541(.A(new_n438), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n589), .ZN(new_n729));
  INV_X1    g543(.A(new_n693), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n269), .B1(new_n261), .B2(new_n278), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n271), .A2(new_n299), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n315), .B1(new_n732), .B2(new_n268), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n291), .A2(new_n292), .A3(new_n734), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n725), .A2(new_n729), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n722), .A2(new_n724), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT106), .B(G143), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G45));
  AOI211_X1 g553(.A(new_n713), .B(new_n660), .C1(new_n396), .C2(new_n399), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n694), .A2(new_n318), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  INV_X1    g556(.A(new_n645), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n663), .B1(new_n725), .B2(new_n659), .ZN(new_n744));
  AOI211_X1 g558(.A(KEYINPUT99), .B(new_n660), .C1(new_n396), .C2(new_n399), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n573), .A2(new_n315), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n573), .A2(new_n749), .A3(new_n315), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(G469), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n586), .A3(new_n668), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(new_n668), .A3(new_n754), .A4(new_n586), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n318), .A2(new_n507), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT41), .B(G113), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  AOI21_X1  g573(.A(new_n682), .B1(new_n679), .B2(new_n395), .ZN(new_n760));
  INV_X1    g574(.A(new_n395), .ZN(new_n761));
  AOI211_X1 g575(.A(KEYINPUT101), .B(new_n761), .C1(new_n676), .C2(new_n678), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n709), .B(new_n686), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n756), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n243), .ZN(G18));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n317), .A2(new_n292), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n450), .B1(new_n767), .B2(new_n701), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n586), .A2(new_n751), .A3(new_n668), .A4(new_n640), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n693), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n730), .A2(new_n752), .A3(new_n641), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(KEYINPUT109), .A3(new_n318), .A4(new_n450), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G119), .ZN(G21));
  NAND2_X1  g589(.A1(new_n438), .A2(new_n640), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n396), .B2(new_n399), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n753), .A2(new_n685), .A3(new_n755), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n301), .A2(new_n269), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n274), .A2(new_n286), .A3(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n666), .A2(G472), .B1(new_n288), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n507), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(G122), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G24));
  NAND4_X1  g599(.A1(new_n740), .A2(new_n693), .A3(new_n769), .A4(new_n781), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G125), .ZN(G27));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n292), .B(new_n317), .C1(new_n701), .C2(new_n788), .ZN(new_n789));
  AOI211_X1 g603(.A(KEYINPUT112), .B(KEYINPUT32), .C1(new_n287), .C2(new_n288), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n507), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n637), .A2(new_n588), .A3(new_n639), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n637), .A2(KEYINPUT111), .A3(new_n588), .A4(new_n639), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n585), .A3(new_n587), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n725), .A2(new_n659), .A3(new_n714), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n794), .A2(new_n795), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n670), .A2(new_n801), .A3(KEYINPUT42), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n700), .A2(new_n705), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n291), .A2(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n701), .A2(new_n788), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(new_n807), .A3(new_n808), .A4(new_n507), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT42), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n318), .A2(new_n740), .A3(new_n507), .A4(new_n797), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n799), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n207), .ZN(G33));
  NAND2_X1  g627(.A1(new_n670), .A2(new_n801), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n706), .A2(new_n506), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n684), .A2(new_n714), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G134), .ZN(G36));
  OR2_X1    g631(.A1(new_n667), .A2(new_n730), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n650), .A2(new_n659), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT43), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT44), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(KEYINPUT44), .A3(new_n823), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n508), .A2(new_n315), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n541), .B1(new_n572), .B2(new_n570), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(KEYINPUT45), .C1(new_n543), .C2(new_n569), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n829), .B1(new_n543), .B2(new_n569), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT45), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n508), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n828), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT46), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n668), .B1(new_n836), .B2(KEYINPUT46), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n586), .B(new_n717), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n826), .A2(new_n801), .A3(new_n827), .A4(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G137), .ZN(G39));
  OAI21_X1  g656(.A(new_n586), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT47), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT47), .B(new_n586), .C1(new_n837), .C2(new_n838), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n318), .A2(new_n800), .A3(new_n507), .A4(new_n796), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  AND2_X1   g664(.A1(new_n751), .A2(new_n668), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n727), .A2(new_n586), .A3(new_n588), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n821), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n735), .A2(new_n506), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n438), .A2(new_n646), .A3(new_n713), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n670), .A2(new_n801), .A3(new_n693), .A4(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n318), .C1(new_n762), .C2(new_n760), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n800), .A2(new_n814), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n781), .A2(new_n693), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n709), .B(new_n714), .C1(new_n760), .C2(new_n762), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n318), .A2(new_n507), .A3(new_n797), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n862), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n667), .A2(new_n507), .A3(new_n670), .A4(new_n686), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n396), .A2(new_n399), .A3(new_n438), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n662), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n695), .B(new_n643), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n799), .A2(new_n809), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n811), .A2(new_n810), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n746), .A2(new_n756), .B1(new_n782), .B2(new_n778), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n764), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(new_n876), .A3(new_n774), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n694), .A2(new_n318), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n866), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n713), .B(KEYINPUT116), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n585), .A2(new_n587), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n735), .A2(new_n730), .A3(new_n777), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n741), .A2(new_n885), .A3(new_n786), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n741), .A2(new_n885), .A3(new_n786), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT52), .B1(new_n888), .B2(new_n715), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n859), .B1(new_n879), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n642), .A2(new_n507), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n666), .A2(G472), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n650), .A2(new_n894), .A3(new_n289), .A4(new_n449), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n768), .A2(new_n893), .B1(new_n895), .B2(new_n707), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n869), .A2(new_n871), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n670), .A2(new_n801), .A3(new_n693), .A4(new_n860), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n706), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n699), .A2(new_n900), .B1(new_n864), .B2(new_n863), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n816), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n812), .ZN(new_n903));
  INV_X1    g717(.A(new_n877), .ZN(new_n904));
  INV_X1    g718(.A(new_n756), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n684), .A3(new_n686), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n904), .A2(new_n906), .A3(new_n774), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n882), .B1(new_n881), .B2(new_n886), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n888), .A2(KEYINPUT52), .A3(new_n715), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(new_n907), .A3(new_n910), .A4(KEYINPUT53), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n892), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n821), .B(KEYINPUT43), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n913), .A2(new_n710), .A3(new_n782), .A4(new_n796), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n851), .A2(new_n587), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n847), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n752), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n801), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n918), .A2(new_n735), .A3(new_n446), .A4(new_n506), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n725), .A2(new_n659), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n919), .A2(KEYINPUT118), .A3(new_n920), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n913), .A2(new_n710), .A3(new_n918), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n864), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n710), .ZN(new_n927));
  INV_X1    g741(.A(new_n782), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n917), .A2(new_n589), .A3(new_n727), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(KEYINPUT50), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n710), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n823), .A2(new_n929), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT50), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n916), .A2(new_n926), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT51), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n916), .A2(new_n926), .A3(new_n935), .A4(KEYINPUT51), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n927), .A2(new_n769), .A3(new_n928), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n919), .B1(new_n744), .B2(new_n745), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n444), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n791), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n925), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT48), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(KEYINPUT48), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n938), .A2(new_n939), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT117), .B1(new_n949), .B2(new_n859), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n891), .A2(new_n911), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(KEYINPUT117), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n912), .B(new_n948), .C1(new_n952), .C2(new_n892), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT119), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT117), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n891), .B2(new_n911), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n957), .B2(new_n950), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(KEYINPUT119), .A3(new_n912), .A4(new_n948), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n443), .A2(new_n264), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT120), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n858), .B1(new_n955), .B2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n264), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n315), .B1(new_n891), .B2(new_n911), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(G210), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n606), .A2(new_n621), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n620), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n965), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n904), .A2(new_n906), .A3(new_n774), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n972), .A2(new_n902), .A3(new_n812), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT53), .B1(new_n973), .B2(new_n910), .ZN(new_n974));
  AND4_X1   g788(.A1(KEYINPUT53), .A2(new_n903), .A3(new_n910), .A4(new_n907), .ZN(new_n975));
  OAI21_X1  g789(.A(G902), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT121), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT121), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n966), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n591), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT56), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n970), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(new_n980), .B2(new_n982), .ZN(G51));
  AND2_X1   g797(.A1(new_n832), .A2(new_n835), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n977), .A2(new_n984), .A3(new_n979), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n828), .B(KEYINPUT57), .ZN(new_n986));
  INV_X1    g800(.A(new_n912), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n892), .B1(new_n891), .B2(new_n911), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n985), .A2(KEYINPUT122), .B1(new_n573), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n977), .A2(new_n991), .A3(new_n984), .A4(new_n979), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n964), .B1(new_n990), .B2(new_n992), .ZN(G54));
  NAND2_X1  g807(.A1(KEYINPUT58), .A2(G475), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n977), .A2(new_n979), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n964), .B1(new_n996), .B2(new_n378), .ZN(new_n997));
  INV_X1    g811(.A(new_n378), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n977), .A2(new_n998), .A3(new_n979), .A4(new_n995), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(G60));
  OAI21_X1  g814(.A(new_n654), .B1(new_n656), .B2(new_n653), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G478), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT59), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1002), .B(new_n1004), .C1(new_n987), .C2(new_n988), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n965), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n958), .A2(new_n912), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1004), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1006), .B1(new_n1008), .B2(new_n1001), .ZN(G63));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT60), .Z(new_n1011));
  NAND3_X1  g825(.A1(new_n951), .A2(new_n691), .A3(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n951), .A2(new_n1011), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n965), .B(new_n1012), .C1(new_n1013), .C2(new_n503), .ZN(new_n1014));
  XNOR2_X1  g828(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G66));
  OAI21_X1  g830(.A(G953), .B1(new_n440), .B2(new_n613), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT124), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n972), .A2(new_n872), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n968), .B1(G898), .B2(new_n264), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G69));
  NAND2_X1  g836(.A1(new_n238), .A2(new_n260), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT125), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(new_n368), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n711), .B2(new_n264), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n841), .A2(new_n876), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n715), .A2(new_n741), .A3(new_n786), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n840), .A2(new_n777), .A3(new_n943), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n849), .A2(new_n1029), .A3(new_n816), .A4(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1026), .B1(new_n1032), .B2(new_n264), .ZN(new_n1033));
  INV_X1    g847(.A(new_n737), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n1034), .A2(KEYINPUT62), .A3(new_n1028), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT62), .B1(new_n1034), .B2(new_n1028), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n318), .A2(new_n507), .ZN(new_n1037));
  NOR4_X1   g851(.A1(new_n723), .A2(new_n1037), .A3(new_n796), .A4(new_n871), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n847), .B2(new_n848), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1035), .A2(new_n841), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1025), .B1(new_n1040), .B2(new_n264), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(G953), .B1(new_n539), .B2(new_n711), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(G72));
  AND3_X1   g858(.A1(new_n261), .A2(new_n278), .A3(new_n269), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1019), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n1027), .A2(new_n1031), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g861(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n702), .A2(new_n315), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1048), .B(new_n1049), .Z(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1045), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1052), .A2(new_n965), .ZN(new_n1053));
  NOR3_X1   g867(.A1(new_n1045), .A2(new_n731), .A3(new_n1051), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n957), .B2(new_n950), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1050), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(new_n731), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(KEYINPUT127), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1057), .A2(new_n1052), .A3(new_n965), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1055), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1058), .A2(new_n1062), .ZN(G57));
endmodule


