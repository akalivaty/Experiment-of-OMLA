

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598;

  XOR2_X1 U327 ( .A(n433), .B(n432), .Z(n295) );
  XOR2_X1 U328 ( .A(n476), .B(KEYINPUT65), .Z(n296) );
  XOR2_X1 U329 ( .A(KEYINPUT40), .B(n508), .Z(n297) );
  XOR2_X1 U330 ( .A(G50GAT), .B(G162GAT), .Z(n429) );
  INV_X1 U331 ( .A(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U332 ( .A(n429), .B(n323), .ZN(n325) );
  XNOR2_X1 U333 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U334 ( .A(n325), .B(n379), .ZN(n326) );
  XNOR2_X1 U335 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U336 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n399) );
  NOR2_X1 U337 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U338 ( .A(n400), .B(n399), .ZN(n574) );
  XNOR2_X1 U339 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U340 ( .A(KEYINPUT36), .ZN(n335) );
  XOR2_X1 U341 ( .A(n333), .B(n332), .Z(n559) );
  XNOR2_X1 U342 ( .A(n497), .B(n496), .ZN(n522) );
  XNOR2_X1 U343 ( .A(n543), .B(n335), .ZN(n596) );
  XNOR2_X1 U344 ( .A(n382), .B(KEYINPUT120), .ZN(n462) );
  XNOR2_X1 U345 ( .A(n463), .B(n462), .ZN(G1350GAT) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U347 ( .A(G1GAT), .B(G183GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n301) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n313) );
  XOR2_X1 U353 ( .A(G57GAT), .B(KEYINPUT13), .Z(n345) );
  XOR2_X1 U354 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U355 ( .A(n345), .B(n428), .Z(n305) );
  XNOR2_X1 U356 ( .A(G78GAT), .B(G211GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U358 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n307) );
  NAND2_X1 U359 ( .A1(G231GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(n309), .B(n308), .Z(n311) );
  XOR2_X1 U362 ( .A(G15GAT), .B(G127GAT), .Z(n458) );
  XNOR2_X1 U363 ( .A(n458), .B(KEYINPUT12), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U365 ( .A(n313), .B(n312), .Z(n556) );
  INV_X1 U366 ( .A(n556), .ZN(n589) );
  INV_X1 U367 ( .A(KEYINPUT78), .ZN(n334) );
  XOR2_X1 U368 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n315) );
  XNOR2_X1 U369 ( .A(G134GAT), .B(KEYINPUT75), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U371 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n317) );
  XNOR2_X1 U372 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n328) );
  XOR2_X1 U375 ( .A(KEYINPUT73), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(n322), .ZN(n349) );
  AND2_X1 U379 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(G36GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n324), .B(G218GAT), .ZN(n379) );
  XOR2_X1 U382 ( .A(n349), .B(n326), .Z(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n330) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G29GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(KEYINPUT69), .B(n331), .ZN(n362) );
  INV_X1 U388 ( .A(n362), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n334), .B(n559), .ZN(n569) );
  INV_X1 U390 ( .A(n569), .ZN(n543) );
  NOR2_X1 U391 ( .A1(n589), .A2(n596), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n336), .B(KEYINPUT45), .ZN(n368) );
  XNOR2_X1 U393 ( .A(G176GAT), .B(G64GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(KEYINPUT74), .ZN(n380) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XNOR2_X1 U396 ( .A(n380), .B(n446), .ZN(n339) );
  AND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n340), .B(KEYINPUT33), .Z(n344) );
  XOR2_X1 U400 ( .A(G78GAT), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n425) );
  XNOR2_X1 U403 ( .A(n425), .B(KEYINPUT32), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U405 ( .A(n346), .B(n345), .Z(n348) );
  XNOR2_X1 U406 ( .A(KEYINPUT31), .B(KEYINPUT71), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n585) );
  XOR2_X1 U409 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n352) );
  XNOR2_X1 U410 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G22GAT), .Z(n354) );
  XNOR2_X1 U413 ( .A(G197GAT), .B(G141GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U415 ( .A(n355), .B(G50GAT), .Z(n357) );
  XOR2_X1 U416 ( .A(G169GAT), .B(G8GAT), .Z(n394) );
  XNOR2_X1 U417 ( .A(n394), .B(G36GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U419 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n359) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n361), .B(n360), .Z(n364) );
  XOR2_X1 U423 ( .A(G113GAT), .B(G1GAT), .Z(n401) );
  XOR2_X1 U424 ( .A(n362), .B(n401), .Z(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n549) );
  INV_X1 U427 ( .A(n549), .ZN(n579) );
  AND2_X1 U428 ( .A1(n585), .A2(n579), .ZN(n367) );
  AND2_X1 U429 ( .A1(n368), .A2(n367), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n369), .B(KEYINPUT109), .ZN(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT41), .B(n585), .ZN(n564) );
  NAND2_X1 U432 ( .A1(n564), .A2(n549), .ZN(n371) );
  XNOR2_X1 U433 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n373) );
  NOR2_X1 U435 ( .A1(n559), .A2(n556), .ZN(n372) );
  AND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n374), .B(KEYINPUT47), .ZN(n375) );
  NAND2_X1 U438 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U439 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n532) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n390) );
  INV_X1 U442 ( .A(KEYINPUT19), .ZN(n381) );
  NAND2_X1 U443 ( .A1(G183GAT), .A2(n381), .ZN(n384) );
  INV_X1 U444 ( .A(G183GAT), .ZN(n382) );
  NAND2_X1 U445 ( .A1(n382), .A2(KEYINPUT19), .ZN(n383) );
  NAND2_X1 U446 ( .A1(n384), .A2(n383), .ZN(n386) );
  XNOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n444) );
  XOR2_X1 U449 ( .A(G211GAT), .B(KEYINPUT86), .Z(n388) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n435) );
  XNOR2_X1 U452 ( .A(n444), .B(n435), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT79), .Z(n392) );
  XNOR2_X1 U455 ( .A(G204GAT), .B(G92GAT), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U457 ( .A(n394), .B(n393), .Z(n396) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n505) );
  INV_X1 U461 ( .A(n505), .ZN(n524) );
  NAND2_X1 U462 ( .A1(n532), .A2(n524), .ZN(n400) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G148GAT), .Z(n403) );
  XOR2_X1 U464 ( .A(G134GAT), .B(KEYINPUT0), .Z(n445) );
  XNOR2_X1 U465 ( .A(n401), .B(n445), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U467 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n405) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n424) );
  XOR2_X1 U470 ( .A(n424), .B(G57GAT), .Z(n407) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n409), .B(n408), .Z(n411) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G162GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(G155GAT), .Z(n413) );
  XNOR2_X1 U477 ( .A(G127GAT), .B(G120GAT), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U479 ( .A(n415), .B(n414), .Z(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U483 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U487 ( .A(n423), .B(n422), .Z(n501) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U489 ( .A(KEYINPUT84), .B(KEYINPUT88), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U492 ( .A(G106GAT), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n295), .B(n434), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n435), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n476) );
  NAND2_X1 U499 ( .A1(n501), .A2(n476), .ZN(n442) );
  OR2_X1 U500 ( .A1(n574), .A2(n442), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n443), .B(KEYINPUT55), .ZN(n461) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U504 ( .A(G113GAT), .B(G176GAT), .Z(n449) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n453) );
  XNOR2_X1 U509 ( .A(G99GAT), .B(KEYINPUT82), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U511 ( .A(G169GAT), .B(n454), .Z(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U513 ( .A(n458), .B(n457), .Z(n460) );
  XNOR2_X1 U514 ( .A(G43GAT), .B(G190GAT), .ZN(n459) );
  XOR2_X1 U515 ( .A(n460), .B(n459), .Z(n507) );
  INV_X1 U516 ( .A(n507), .ZN(n535) );
  NAND2_X1 U517 ( .A1(n461), .A2(n535), .ZN(n570) );
  NOR2_X1 U518 ( .A1(n589), .A2(n570), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n579), .A2(n570), .ZN(n465) );
  XNOR2_X1 U520 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(G1348GAT) );
  NAND2_X1 U522 ( .A1(n585), .A2(n549), .ZN(n498) );
  NOR2_X1 U523 ( .A1(n589), .A2(n543), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT16), .ZN(n481) );
  NOR2_X1 U525 ( .A1(n535), .A2(n476), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT95), .ZN(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT26), .B(n468), .ZN(n576) );
  XNOR2_X1 U528 ( .A(n505), .B(KEYINPUT27), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n576), .A2(n475), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n524), .A2(n535), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n476), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT96), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n474) );
  INV_X1 U535 ( .A(n501), .ZN(n575) );
  NOR2_X1 U536 ( .A1(n474), .A2(n575), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n475), .A2(n501), .ZN(n533) );
  XOR2_X1 U538 ( .A(KEYINPUT28), .B(n296), .Z(n529) );
  INV_X1 U539 ( .A(n529), .ZN(n534) );
  NAND2_X1 U540 ( .A1(n533), .A2(n534), .ZN(n477) );
  NOR2_X1 U541 ( .A1(n535), .A2(n477), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n480), .B(KEYINPUT97), .ZN(n493) );
  NAND2_X1 U543 ( .A1(n481), .A2(n493), .ZN(n511) );
  NOR2_X1 U544 ( .A1(n498), .A2(n511), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n488), .A2(n575), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n488), .A2(n524), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n484), .B(KEYINPUT98), .ZN(n485) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(n485), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U552 ( .A1(n488), .A2(n535), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n490) );
  NAND2_X1 U555 ( .A1(n488), .A2(n529), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n596), .A2(n556), .ZN(n492) );
  NAND2_X1 U559 ( .A1(n493), .A2(n492), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n495) );
  INV_X1 U561 ( .A(KEYINPUT101), .ZN(n494) );
  NOR2_X1 U562 ( .A1(n522), .A2(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n509), .A2(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n509), .A2(n505), .ZN(n506) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n507), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n297), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n509), .A2(n534), .ZN(n510) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  NAND2_X1 U576 ( .A1(n579), .A2(n564), .ZN(n521) );
  NOR2_X1 U577 ( .A1(n521), .A2(n511), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n575), .A2(n517), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n524), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U582 ( .A(G71GAT), .B(KEYINPUT105), .Z(n516) );
  NAND2_X1 U583 ( .A1(n517), .A2(n535), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n519) );
  NAND2_X1 U586 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n575), .A2(n528), .ZN(n523) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U595 ( .A1(n528), .A2(n535), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n548), .A2(n536), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n549), .A2(n544), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U606 ( .A1(n544), .A2(n564), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT111), .B(KEYINPUT50), .Z(n541) );
  NAND2_X1 U609 ( .A1(n544), .A2(n556), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n576), .A2(n548), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT114), .Z(n552) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT113), .B(n553), .Z(n555) );
  NAND2_X1 U623 ( .A1(n560), .A2(n564), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U626 ( .A1(n560), .A2(n556), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n562) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  INV_X1 U632 ( .A(n564), .ZN(n565) );
  NOR2_X1 U633 ( .A1(n565), .A2(n570), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n568), .ZN(G1349GAT) );
  INV_X1 U637 ( .A(KEYINPUT58), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(G190GAT), .ZN(G1351GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n578) );
  INV_X1 U642 ( .A(n576), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n595) );
  NOR2_X1 U644 ( .A1(n579), .A2(n595), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT121), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT59), .B(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n595), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT61), .B(KEYINPUT123), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(G204GAT), .B(n588), .Z(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n595), .ZN(n591) );
  XNOR2_X1 U655 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(G211GAT), .B(n592), .ZN(G1354GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n594) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(n598) );
  NOR2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U662 ( .A(n598), .B(n597), .Z(G1355GAT) );
endmodule

