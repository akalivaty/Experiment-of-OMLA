//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n451), .B2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT70), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT71), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n470), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(new_n471), .B1(new_n472), .B2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT72), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n470), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n469), .A2(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n470), .A2(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n478), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G88), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n513), .B2(new_n514), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT74), .B1(new_n520), .B2(new_n511), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT7), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n508), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(G51), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n505), .A2(new_n506), .ZN(new_n528));
  INV_X1    g103(.A(new_n502), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n531), .A2(G90), .B1(G52), .B2(new_n526), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n519), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT76), .B(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n531), .A2(new_n545), .B1(G43), .B2(new_n526), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n528), .A2(new_n529), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n525), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n508), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n530), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n508), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n568), .A2(KEYINPUT79), .A3(G91), .A4(new_n569), .ZN(new_n573));
  AOI211_X1 g148(.A(new_n554), .B(new_n565), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  INV_X1    g150(.A(new_n565), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT80), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n526), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n568), .A2(G87), .A3(new_n569), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(KEYINPUT81), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n568), .A2(new_n585), .A3(G87), .A4(new_n569), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n526), .A2(G48), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n519), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n568), .A2(G86), .A3(new_n569), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT82), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n568), .A2(new_n593), .A3(G86), .A4(new_n569), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n519), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n530), .A2(new_n599), .B1(new_n600), .B2(new_n525), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  OR3_X1    g179(.A1(G171), .A2(KEYINPUT83), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT83), .B1(G171), .B2(new_n604), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT85), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n570), .B2(new_n609), .ZN(new_n610));
  AND4_X1   g185(.A1(KEYINPUT78), .A2(new_n528), .A3(new_n529), .A4(new_n508), .ZN(new_n611));
  AOI21_X1  g186(.A(KEYINPUT78), .B1(new_n507), .B2(new_n508), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n608), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n613), .A2(G92), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n556), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n605), .B(new_n606), .C1(G868), .C2(new_n622), .ZN(G284));
  OAI211_X1 g198(.A(new_n605), .B(new_n606), .C1(G868), .C2(new_n622), .ZN(G321));
  NAND2_X1  g199(.A1(G168), .A2(G868), .ZN(new_n625));
  XOR2_X1   g200(.A(G299), .B(KEYINPUT86), .Z(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT87), .Z(G297));
  XOR2_X1   g203(.A(new_n627), .B(KEYINPUT88), .Z(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n622), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n544), .A2(new_n546), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n604), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n621), .A2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n469), .A2(new_n472), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT91), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n482), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n484), .A2(G123), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT92), .B(G2096), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n640), .A2(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT90), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n642), .A2(new_n649), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT94), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G2451), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(KEYINPUT94), .ZN(new_n664));
  INV_X1    g239(.A(G2451), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(new_n663), .B2(new_n666), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n659), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n662), .A2(G2451), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g250(.A1(new_n675), .A2(new_n656), .A3(new_n658), .A4(new_n669), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT93), .B(KEYINPUT16), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G2454), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G14), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n678), .B1(new_n672), .B2(new_n676), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT95), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT95), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n683), .A2(new_n684), .A3(G14), .A4(new_n679), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G401));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT96), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2072), .B(G2078), .Z(new_n691));
  XNOR2_X1  g266(.A(G2084), .B(G2090), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT18), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT97), .B(KEYINPUT17), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n692), .C1(new_n697), .C2(new_n690), .ZN(new_n698));
  INV_X1    g273(.A(new_n692), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n690), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n694), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G2096), .B(G2100), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(G227));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1971), .B(G1976), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT19), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1956), .B(G2474), .Z(new_n711));
  XOR2_X1   g286(.A(G1961), .B(G1966), .Z(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(new_n713), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT20), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT98), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(KEYINPUT98), .B1(new_n717), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n707), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT99), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n717), .A2(new_n719), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT98), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n729), .A2(new_n720), .A3(new_n706), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n723), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n723), .B2(new_n730), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n705), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n733), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n735), .A2(new_n704), .A3(new_n731), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(G229));
  NAND2_X1  g312(.A1(new_n622), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G4), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1348), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NOR2_X1   g317(.A1(G162), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G35), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT106), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT29), .Z(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G2090), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(KEYINPUT107), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(KEYINPUT107), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(G299), .A2(G16), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1956), .Z(new_n756));
  INV_X1    g331(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n747), .A2(G2090), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n470), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT103), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n482), .A2(G139), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n769));
  OAI21_X1  g344(.A(G29), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G33), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(G29), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G2072), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n752), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n752), .B2(G19), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G1341), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n752), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n752), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1966), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(KEYINPUT24), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT24), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n474), .B2(new_n742), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT104), .ZN(new_n788));
  INV_X1    g363(.A(new_n647), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n789), .A2(G29), .B1(new_n786), .B2(new_n785), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n742), .A2(G27), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n499), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2078), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G28), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n742), .B1(new_n795), .B2(G28), .ZN(new_n797));
  AND2_X1   g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NOR2_X1   g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n792), .B2(new_n793), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n788), .A2(new_n790), .A3(new_n794), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n787), .A2(KEYINPUT104), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n781), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT105), .B1(new_n772), .B2(G2072), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n772), .A2(KEYINPUT105), .A3(G2072), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n778), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G128), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(new_n481), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n809), .A2(G140), .A3(new_n470), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(G116), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT102), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n742), .A2(G26), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT28), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n740), .B2(new_n739), .ZN(new_n823));
  NOR2_X1   g398(.A1(G171), .A2(new_n752), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G5), .B2(new_n752), .ZN(new_n825));
  INV_X1    g400(.A(G1961), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n482), .A2(G141), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n484), .A2(G129), .ZN(new_n830));
  NAND3_X1  g405(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT26), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n833), .A2(new_n834), .B1(G105), .B2(new_n472), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n829), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G29), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n742), .A2(G32), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT27), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(KEYINPUT27), .ZN(new_n841));
  INV_X1    g416(.A(G1996), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n827), .A2(new_n828), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n807), .A2(new_n823), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n750), .A2(new_n759), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT109), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n750), .A2(new_n759), .A3(new_n846), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT109), .B1(new_n852), .B2(new_n849), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(G107), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(G2105), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n484), .B2(G119), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n482), .A2(G131), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  MUX2_X1   g434(.A(G25), .B(new_n859), .S(G29), .Z(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G1991), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT100), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n860), .B(new_n862), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n752), .A2(G24), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n602), .B2(new_n752), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(G1986), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n752), .A2(G23), .ZN(new_n868));
  INV_X1    g443(.A(G288), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n752), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT33), .B(G1976), .Z(new_n871));
  XOR2_X1   g446(.A(new_n870), .B(new_n871), .Z(new_n872));
  NOR2_X1   g447(.A1(G16), .A2(G22), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G166), .B2(G16), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(G1971), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n752), .A2(G6), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n595), .B2(new_n752), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT32), .B(G1981), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT34), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n867), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(KEYINPUT34), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT36), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(KEYINPUT36), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n851), .A2(new_n853), .B1(new_n891), .B2(new_n892), .ZN(G311));
  INV_X1    g468(.A(new_n890), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n889), .B1(new_n883), .B2(new_n884), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n852), .A2(KEYINPUT109), .A3(new_n849), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G150));
  AOI22_X1  g474(.A1(new_n531), .A2(G93), .B1(G55), .B2(new_n526), .ZN(new_n900));
  NAND2_X1  g475(.A1(G80), .A2(G543), .ZN(new_n901));
  INV_X1    g476(.A(G67), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n556), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G651), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT110), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT111), .B(G860), .Z(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT112), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT37), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n547), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n632), .A2(new_n905), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n622), .A2(G559), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT39), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n913), .B1(new_n920), .B2(new_n910), .ZN(G145));
  NAND2_X1  g496(.A1(new_n815), .A2(new_n499), .ZN(new_n922));
  NAND4_X1  g497(.A1(G164), .A2(new_n808), .A3(new_n810), .A4(new_n814), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n769), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n767), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n922), .B(new_n923), .C1(new_n768), .C2(new_n769), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n836), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n482), .A2(G142), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n484), .A2(G130), .ZN(new_n931));
  OR2_X1    g506(.A1(G106), .A2(G2105), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n932), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n857), .A2(KEYINPUT113), .A3(new_n858), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT113), .B1(new_n857), .B2(new_n858), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n638), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n859), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n638), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n935), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n943), .A3(new_n935), .ZN(new_n946));
  INV_X1    g521(.A(new_n836), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n926), .A2(new_n927), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n929), .A2(new_n945), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n926), .A2(new_n927), .A3(new_n947), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n947), .B1(new_n926), .B2(new_n927), .ZN(new_n951));
  INV_X1    g526(.A(new_n946), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n950), .A2(new_n951), .B1(new_n952), .B2(new_n944), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n647), .B(G160), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(G162), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(KEYINPUT114), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n952), .A2(new_n944), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n948), .A4(new_n929), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n955), .B(G162), .Z(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n961), .A3(new_n953), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g540(.A(new_n916), .B(new_n634), .Z(new_n966));
  NAND2_X1  g541(.A1(new_n575), .A2(new_n576), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n554), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n575), .A2(KEYINPUT80), .A3(new_n576), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n622), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n621), .B1(new_n574), .B2(new_n577), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT41), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT41), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n916), .B(new_n634), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(KEYINPUT115), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT115), .B1(new_n974), .B2(new_n977), .ZN(new_n979));
  XNOR2_X1  g554(.A(G288), .B(new_n595), .ZN(new_n980));
  XNOR2_X1  g555(.A(G166), .B(new_n602), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n978), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n982), .B(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(KEYINPUT115), .A3(new_n977), .A4(new_n974), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G868), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(new_n909), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G868), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n604), .B1(new_n984), .B2(new_n987), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT116), .B1(new_n995), .B2(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(G295));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n993), .ZN(G331));
  NAND2_X1  g573(.A1(G171), .A2(G286), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G171), .A2(G286), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(new_n914), .B2(new_n915), .ZN(new_n1002));
  XNOR2_X1  g577(.A(G301), .B(G286), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n916), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT41), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n976), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT41), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n976), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n982), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G37), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n972), .B2(new_n973), .ZN(new_n1015));
  INV_X1    g590(.A(new_n982), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1010), .ZN(new_n1020));
  AOI21_X1  g595(.A(G37), .B1(new_n1020), .B2(new_n982), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1017), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1024), .B(new_n1025), .ZN(G397));
  INV_X1    g601(.A(KEYINPUT126), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n836), .B(new_n842), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n815), .B(new_n821), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n499), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n468), .A2(G40), .A3(new_n473), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n859), .A2(new_n862), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n859), .A2(new_n862), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1038), .B(new_n1040), .C1(new_n1035), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n602), .B(G1986), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1036), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n499), .A2(new_n1031), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1033), .B1(new_n1050), .B2(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n499), .A2(new_n1053), .A3(new_n1031), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1033), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1971), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n518), .A2(new_n521), .A3(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n518), .A2(new_n521), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1060), .B(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1050), .A2(new_n1033), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  INV_X1    g646(.A(new_n590), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n593), .B1(new_n613), .B2(G86), .ZN(new_n1073));
  INV_X1    g648(.A(new_n594), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1071), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n531), .A2(G86), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G1981), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1070), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n583), .A2(KEYINPUT81), .ZN(new_n1083));
  INV_X1    g658(.A(new_n582), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(G1976), .A3(new_n586), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n584), .A2(KEYINPUT118), .A3(G1976), .A4(new_n586), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1069), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1081), .A2(new_n1082), .B1(KEYINPUT52), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1976), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(G288), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(new_n1087), .A3(new_n1069), .A4(new_n1088), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1066), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1058), .A3(new_n1034), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1098), .B2(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1050), .A2(KEYINPUT50), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n1034), .A3(new_n1054), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n826), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1057), .A2(KEYINPUT53), .A3(new_n793), .A4(new_n1058), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1099), .A2(G301), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1100), .A2(new_n786), .A3(new_n1034), .A4(new_n1054), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1111), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1112));
  OAI211_X1 g687(.A(G168), .B(new_n1110), .C1(new_n1112), .C2(G1966), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  INV_X1    g689(.A(G1966), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1098), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(G168), .B1(new_n1116), .B2(new_n1110), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1119), .A3(G8), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1105), .A2(KEYINPUT54), .A3(new_n1106), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1109), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n967), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n575), .A2(new_n576), .A3(new_n1124), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT120), .B(G1956), .Z(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1101), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT56), .B(G2072), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1112), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1126), .A2(new_n1127), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1127), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1124), .B1(new_n575), .B2(new_n576), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1348), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1050), .A2(new_n1033), .A3(G2067), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(new_n621), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1140), .A2(KEYINPUT122), .A3(new_n621), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1133), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1126), .A2(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT58), .B(G1341), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1098), .A2(G1996), .B1(new_n1067), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n547), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1154), .A3(new_n547), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1153), .A2(new_n1155), .B1(new_n1140), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n622), .A2(new_n1139), .A3(new_n1138), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT60), .B1(new_n1158), .B2(new_n1141), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1137), .A2(new_n1133), .A3(KEYINPUT61), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1149), .A2(new_n1157), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1123), .B1(new_n1145), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1118), .A2(new_n1163), .A3(new_n1120), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1105), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1113), .A2(new_n1119), .A3(G8), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1110), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1966), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1169));
  OAI21_X1  g744(.A(G286), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(G8), .A3(new_n1113), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1171), .B2(KEYINPUT51), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT123), .B1(new_n1172), .B2(new_n1163), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1121), .A2(new_n1174), .A3(KEYINPUT62), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1166), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1095), .B1(new_n1162), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT119), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1179));
  AOI211_X1 g754(.A(G1981), .B(new_n590), .C1(new_n592), .C2(new_n594), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1071), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1080), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(new_n1069), .A3(new_n1082), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(KEYINPUT119), .A4(new_n1093), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1178), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1183), .A2(new_n1091), .A3(new_n869), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1069), .B1(new_n1188), .B2(new_n1180), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1183), .A2(new_n1184), .A3(new_n1093), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1185), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1068), .B(G286), .C1(new_n1116), .C2(new_n1110), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1195), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1066), .A2(new_n1090), .A3(new_n1093), .A4(new_n1195), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1194), .A2(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1190), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1049), .B1(new_n1177), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1029), .B(new_n947), .C1(new_n1202), .C2(G1996), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1036), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1035), .B2(G1996), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT125), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT47), .ZN(new_n1208));
  NOR3_X1   g783(.A1(G290), .A2(new_n1035), .A3(G1986), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT48), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1208), .B1(new_n1045), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n815), .A2(G2067), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1035), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1215), .A2(KEYINPUT124), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1215), .A2(KEYINPUT124), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1211), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1027), .B1(new_n1201), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1049), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1161), .A2(new_n1145), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1123), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1105), .B1(new_n1172), .B2(new_n1163), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1174), .B1(new_n1121), .B2(KEYINPUT62), .ZN(new_n1226));
  AOI211_X1 g801(.A(KEYINPUT123), .B(new_n1163), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1094), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1195), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1231), .B1(new_n1193), .B2(new_n1185), .ZN(new_n1232));
  OAI211_X1 g807(.A(new_n1187), .B(new_n1189), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1221), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1234), .A2(KEYINPUT126), .A3(new_n1218), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1220), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g811(.A1(G227), .A2(new_n460), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n686), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g813(.A(new_n1239), .B1(new_n734), .B2(new_n736), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n964), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g815(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g816(.A(KEYINPUT127), .B1(new_n1024), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1244));
  AOI211_X1 g818(.A(new_n1244), .B(new_n1241), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1245));
  NOR2_X1   g819(.A1(new_n1243), .A2(new_n1245), .ZN(G308));
  AOI21_X1  g820(.A(new_n1022), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1247));
  AND4_X1   g821(.A1(new_n1022), .A2(new_n1012), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1248));
  OAI21_X1  g822(.A(new_n1242), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g823(.A1(new_n1249), .A2(new_n1244), .ZN(new_n1250));
  NAND3_X1  g824(.A1(new_n1024), .A2(KEYINPUT127), .A3(new_n1242), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n1250), .A2(new_n1251), .ZN(G225));
endmodule


