//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n447, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(KEYINPUT68), .B(new_n462), .C1(new_n463), .C2(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n463), .B2(KEYINPUT68), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G113), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n463), .ZN(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n469), .A2(new_n470), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n469), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR3_X1   g062(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT71), .Z(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n475), .A2(new_n476), .ZN(new_n495));
  AND4_X1   g070(.A1(new_n494), .A2(new_n495), .A3(G138), .A4(new_n470), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n469), .A2(G138), .A3(new_n470), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n469), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n470), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n507), .A2(new_n509), .B1(KEYINPUT5), .B2(new_n506), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(new_n517), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT74), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n517), .A2(new_n506), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G651), .B1(G50), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AND3_X1   g109(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n535));
  AOI211_X1 g110(.A(new_n534), .B(new_n535), .C1(G51), .C2(new_n529), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n523), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n529), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(new_n522), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n513), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n523), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n512), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(G43), .B2(new_n529), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n512), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n529), .A2(G53), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(KEYINPUT76), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n529), .A2(G53), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n518), .A2(G91), .A3(new_n522), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n523), .A2(G87), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n519), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G49), .B2(new_n529), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n523), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n512), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G48), .B2(new_n529), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n579), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n580), .A2(new_n579), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n529), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n513), .B2(new_n590), .C1(new_n541), .C2(new_n591), .ZN(G290));
  AND3_X1   g167(.A1(new_n518), .A2(G92), .A3(new_n522), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n529), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  XNOR2_X1  g178(.A(G321), .B(KEYINPUT79), .ZN(G284));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n573), .B(KEYINPUT80), .Z(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(new_n600), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n484), .B2(G135), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n486), .A2(KEYINPUT81), .A3(G123), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n499), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT84), .Z(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT86), .Z(new_n655));
  OAI21_X1  g230(.A(new_n653), .B1(new_n649), .B2(new_n651), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n650), .B2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n649), .A3(new_n651), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n655), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n670), .A2(KEYINPUT20), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n671), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(new_n667), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n673), .B(new_n675), .C1(KEYINPUT20), .C2(new_n670), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1991), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G35), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G162), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT29), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2090), .ZN(new_n687));
  INV_X1    g262(.A(G1961), .ZN(new_n688));
  NOR2_X1   g263(.A1(G5), .A2(G16), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(G301), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n687), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT95), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT26), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n484), .A2(G141), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n486), .A2(G129), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G29), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n683), .A2(G33), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  AOI22_X1  g287(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  INV_X1    g288(.A(G139), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n712), .B1(new_n713), .B2(new_n470), .C1(new_n483), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n715), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2072), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G28), .ZN(new_n719));
  OR2_X1    g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n719), .A2(new_n683), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n624), .A2(new_n683), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n716), .A2(new_n717), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n718), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n683), .B1(new_n726), .B2(G34), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(new_n726), .B2(G34), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(new_n727), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n481), .B2(new_n683), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n708), .A2(new_n709), .A3(new_n725), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G21), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G168), .B2(G16), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT96), .B(G1966), .Z(new_n737));
  XOR2_X1   g312(.A(new_n736), .B(new_n737), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n731), .A2(new_n732), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT94), .Z(new_n740));
  NOR2_X1   g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n683), .A2(G26), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n744));
  INV_X1    g319(.A(G140), .ZN(new_n745));
  INV_X1    g320(.A(G128), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n744), .B1(new_n483), .B2(new_n745), .C1(new_n746), .C2(new_n499), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n742), .B1(new_n747), .B2(G29), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n742), .B(new_n748), .S(KEYINPUT28), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n691), .A2(G4), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n600), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n734), .A2(new_n741), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n683), .A2(G27), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT99), .Z(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n683), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT100), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT90), .B(G16), .ZN(new_n761));
  INV_X1    g336(.A(G19), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n554), .B2(new_n761), .ZN(new_n764));
  MUX2_X1   g339(.A(new_n763), .B(new_n764), .S(KEYINPUT92), .Z(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  NOR3_X1   g341(.A1(new_n755), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n693), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G20), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  INV_X1    g348(.A(new_n752), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(G1956), .B1(new_n774), .B2(G1348), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n692), .A2(new_n688), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n775), .B1(G1956), .B2(new_n773), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n768), .A2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G22), .B(G303), .S(new_n761), .Z(new_n782));
  INV_X1    g357(.A(G1971), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n691), .B1(new_n586), .B2(new_n587), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT32), .B(G1981), .Z(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n691), .A2(G6), .ZN(new_n788));
  OR3_X1    g363(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n787), .B1(new_n785), .B2(new_n788), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n784), .A2(new_n789), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT91), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(KEYINPUT91), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n797), .A2(KEYINPUT34), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G25), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n484), .A2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n486), .A2(G119), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT88), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT89), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n804), .B1(new_n811), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT35), .B(G1991), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G24), .B(G290), .S(new_n761), .Z(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n803), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n803), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n781), .B1(new_n821), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n823), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n825), .A2(new_n780), .A3(new_n768), .ZN(G150));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n610), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n523), .A2(G93), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n529), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n512), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G651), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(KEYINPUT102), .A3(G651), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n830), .A2(new_n831), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n555), .B(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n829), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n829), .A2(new_n840), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(G164), .B(new_n747), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n715), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n704), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n810), .B(new_n627), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n484), .A2(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n470), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G130), .B2(new_n486), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n850), .B(new_n855), .Z(new_n856));
  AND2_X1   g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n849), .A2(new_n856), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT103), .ZN(new_n859));
  XNOR2_X1  g434(.A(G160), .B(new_n624), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n492), .B(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n858), .B2(KEYINPUT103), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n864), .A2(new_n865), .A3(new_n861), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n864), .B2(new_n861), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g444(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT106), .Z(new_n871));
  XNOR2_X1  g446(.A(G288), .B(G290), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n586), .A2(G303), .A3(new_n587), .ZN(new_n874));
  AOI21_X1  g449(.A(G303), .B1(new_n586), .B2(new_n587), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(G305), .A2(G166), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n586), .A2(G303), .A3(new_n587), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n839), .B(new_n554), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n612), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n594), .A2(G299), .A3(new_n599), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(G299), .B1(new_n594), .B2(new_n599), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n600), .A2(new_n573), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n884), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n882), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n882), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n871), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n871), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n839), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(G868), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(G295));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n909), .A3(new_n907), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n902), .B1(new_n901), .B2(new_n897), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n898), .A2(new_n871), .A3(new_n899), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n601), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n913), .B2(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n544), .A2(G286), .A3(new_n546), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G286), .B1(new_n544), .B2(new_n546), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n918), .A2(new_n840), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G301), .A2(G168), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n883), .B1(new_n921), .B2(new_n917), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n892), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n840), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n883), .A3(new_n917), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n895), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n926), .A3(new_n880), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n880), .A2(KEYINPUT108), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n876), .A2(new_n879), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n930), .B2(new_n934), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT43), .B(new_n929), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n930), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n927), .A2(new_n928), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n916), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n939), .B(new_n929), .C1(new_n936), .C2(new_n937), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n916), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n945), .B2(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT110), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n498), .B2(new_n503), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n471), .A2(G40), .A3(new_n480), .A4(new_n472), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  AND2_X1   g536(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n962));
  NOR2_X1   g537(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n963));
  OAI21_X1  g538(.A(G125), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n478), .B2(new_n463), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n965), .B2(G2105), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n472), .A4(new_n471), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n957), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT46), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(KEYINPUT46), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n747), .B(G2067), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(new_n703), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  INV_X1    g552(.A(new_n968), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n968), .A2(new_n974), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT113), .Z(new_n980));
  NOR2_X1   g555(.A1(new_n704), .A2(new_n969), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n968), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n971), .A2(new_n704), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT112), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(new_n814), .A3(new_n811), .A4(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n747), .A2(G2067), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n984), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n810), .B(new_n813), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n968), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT48), .Z(new_n992));
  AOI211_X1 g567(.A(new_n977), .B(new_n987), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G303), .A2(G8), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT55), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n960), .A2(new_n967), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT45), .B(new_n954), .C1(new_n498), .C2(new_n503), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n957), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n783), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n954), .C1(new_n498), .C2(new_n503), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n997), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(G2090), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n996), .A2(G8), .A3(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1001), .A2(new_n997), .A3(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(new_n999), .B2(new_n783), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n995), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n999), .B2(G2078), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1004), .A2(new_n688), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OR3_X1    g591(.A1(new_n999), .A2(new_n1013), .A3(G2078), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G171), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n580), .A2(new_n1021), .A3(new_n584), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n580), .B2(new_n584), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1024), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n1028));
  INV_X1    g603(.A(new_n496), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n501), .A2(new_n502), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n486), .B2(G126), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1010), .B1(new_n1033), .B2(new_n997), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1027), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n1034), .C1(new_n1036), .C2(G288), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1034), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G288), .A2(new_n1036), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1012), .A2(new_n1019), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1007), .A2(new_n1044), .A3(new_n732), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n999), .A2(new_n737), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT116), .B1(new_n1004), .B2(G2084), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n1010), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(KEYINPUT51), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(G8), .C1(new_n1048), .C2(G286), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1043), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT127), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1043), .A2(KEYINPUT127), .A3(new_n1057), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1023), .B1(new_n1035), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1039), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1069), .B1(new_n1072), .B2(new_n1006), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1049), .A2(G286), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(KEYINPUT63), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1042), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1078), .A3(new_n1076), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1073), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1064), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1013), .B(G2078), .C1(new_n958), .C2(KEYINPUT124), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n958), .A2(KEYINPUT124), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n957), .A2(new_n1085), .A3(new_n998), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1016), .A2(G301), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT54), .B1(new_n1019), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(G301), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1014), .A2(new_n1015), .A3(new_n1087), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1093), .A2(KEYINPUT126), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT126), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1090), .B(new_n1062), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n573), .A2(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n571), .B2(new_n572), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1004), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n957), .A2(new_n997), .A3(new_n998), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1108), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n600), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1033), .A2(new_n997), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  INV_X1    g690(.A(G2067), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1033), .A2(new_n997), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1004), .A2(new_n753), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1115), .A2(new_n1122), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1111), .B1(new_n1113), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n609), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1123), .A2(new_n1121), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n600), .A4(new_n1120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1106), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1108), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(KEYINPUT119), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  AND3_X1   g719(.A1(new_n1033), .A2(new_n997), .A3(new_n1117), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1117), .B1(new_n1033), .B2(new_n997), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n957), .A2(new_n969), .A3(new_n997), .A4(new_n998), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1143), .B1(new_n1149), .B2(new_n555), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1143), .B2(KEYINPUT120), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n554), .B(new_n1152), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1141), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1152), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1149), .A2(new_n555), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n554), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1156), .B(KEYINPUT121), .C1(new_n1157), .C2(new_n1143), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1140), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1132), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(KEYINPUT122), .B(new_n1140), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1125), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1102), .B1(new_n1163), .B2(KEYINPUT123), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1125), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1083), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(G290), .B(G1986), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n990), .B1(new_n978), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n993), .B1(new_n1167), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(G319), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G227), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n647), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G229), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1175), .A2(new_n868), .A3(new_n947), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


