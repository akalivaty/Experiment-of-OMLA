

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781;

  NAND2_X1 U372 ( .A1(n644), .A2(n641), .ZN(n771) );
  XNOR2_X1 U373 ( .A(n604), .B(n603), .ZN(n780) );
  XNOR2_X1 U374 ( .A(n531), .B(KEYINPUT40), .ZN(n673) );
  XNOR2_X1 U375 ( .A(n471), .B(n470), .ZN(n629) );
  INV_X1 U376 ( .A(G902), .ZN(n407) );
  AND2_X1 U377 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X2 U378 ( .A1(n389), .A2(n387), .ZN(n747) );
  BUF_X1 U379 ( .A(n747), .Z(n751) );
  INV_X1 U380 ( .A(G953), .ZN(n772) );
  AND2_X1 U381 ( .A1(n377), .A2(n380), .ZN(n376) );
  AND2_X2 U382 ( .A1(n404), .A2(n402), .ZN(n602) );
  XNOR2_X2 U383 ( .A(G116), .B(G113), .ZN(n459) );
  XNOR2_X2 U384 ( .A(n482), .B(n481), .ZN(n758) );
  XNOR2_X2 U385 ( .A(KEYINPUT65), .B(G143), .ZN(n446) );
  XNOR2_X2 U386 ( .A(n552), .B(n551), .ZN(n589) );
  NOR2_X1 U387 ( .A1(n627), .A2(n597), .ZN(n598) );
  NAND2_X1 U388 ( .A1(n638), .A2(n637), .ZN(n396) );
  NAND2_X1 U389 ( .A1(n385), .A2(n383), .ZN(n382) );
  NOR2_X1 U390 ( .A1(n624), .A2(n623), .ZN(n725) );
  NOR2_X1 U391 ( .A1(n631), .A2(n393), .ZN(n412) );
  XNOR2_X1 U392 ( .A(n598), .B(n599), .ZN(n605) );
  XNOR2_X1 U393 ( .A(n459), .B(n458), .ZN(n461) );
  INV_X1 U394 ( .A(KEYINPUT3), .ZN(n458) );
  XNOR2_X1 U395 ( .A(KEYINPUT18), .B(G125), .ZN(n484) );
  AND2_X1 U396 ( .A1(n682), .A2(n351), .ZN(n388) );
  AND2_X1 U397 ( .A1(n417), .A2(KEYINPUT66), .ZN(n351) );
  XNOR2_X2 U398 ( .A(n371), .B(KEYINPUT79), .ZN(n625) );
  XNOR2_X2 U399 ( .A(n363), .B(n394), .ZN(n644) );
  NAND2_X2 U400 ( .A1(n602), .A2(n696), .ZN(n371) );
  XNOR2_X2 U401 ( .A(n457), .B(n456), .ZN(n393) );
  XNOR2_X2 U402 ( .A(n494), .B(n493), .ZN(n550) );
  XNOR2_X2 U403 ( .A(n583), .B(KEYINPUT33), .ZN(n686) );
  XNOR2_X2 U404 ( .A(n488), .B(n448), .ZN(n467) );
  NAND2_X1 U405 ( .A1(n408), .A2(n407), .ZN(n406) );
  INV_X1 U406 ( .A(G469), .ZN(n408) );
  NAND2_X1 U407 ( .A1(G902), .A2(G469), .ZN(n410) );
  AND2_X1 U408 ( .A1(n536), .A2(n547), .ZN(n554) );
  NOR2_X1 U409 ( .A1(n541), .A2(n629), .ZN(n535) );
  INV_X1 U410 ( .A(n406), .ZN(n400) );
  AND2_X1 U411 ( .A1(G953), .A2(G902), .ZN(n476) );
  INV_X1 U412 ( .A(G128), .ZN(n445) );
  INV_X1 U413 ( .A(KEYINPUT86), .ZN(n394) );
  NOR2_X1 U414 ( .A1(n622), .A2(n533), .ZN(n534) );
  XNOR2_X1 U415 ( .A(G104), .B(G110), .ZN(n450) );
  XNOR2_X1 U416 ( .A(KEYINPUT16), .B(G122), .ZN(n481) );
  XNOR2_X1 U417 ( .A(n431), .B(n366), .ZN(n521) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U420 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U421 ( .A(n522), .B(KEYINPUT105), .ZN(n367) );
  AND2_X1 U422 ( .A1(n379), .A2(n378), .ZN(n374) );
  INV_X1 U423 ( .A(KEYINPUT19), .ZN(n551) );
  NAND2_X1 U424 ( .A1(n550), .A2(n549), .ZN(n552) );
  OR2_X1 U425 ( .A1(n674), .A2(G902), .ZN(n471) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n506) );
  XNOR2_X1 U427 ( .A(n420), .B(n435), .ZN(n440) );
  NAND2_X1 U428 ( .A1(n646), .A2(G234), .ZN(n420) );
  NAND2_X1 U429 ( .A1(n400), .A2(n546), .ZN(n399) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n492) );
  XNOR2_X1 U431 ( .A(G134), .B(G131), .ZN(n447) );
  XNOR2_X1 U432 ( .A(KEYINPUT69), .B(G101), .ZN(n464) );
  INV_X1 U433 ( .A(KEYINPUT72), .ZN(n424) );
  XOR2_X1 U434 ( .A(KEYINPUT106), .B(KEYINPUT104), .Z(n515) );
  XNOR2_X1 U435 ( .A(G134), .B(G122), .ZN(n514) );
  XNOR2_X1 U436 ( .A(G116), .B(G107), .ZN(n517) );
  XOR2_X1 U437 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n508) );
  XNOR2_X1 U438 ( .A(G113), .B(G131), .ZN(n500) );
  XOR2_X1 U439 ( .A(G104), .B(G143), .Z(n501) );
  XNOR2_X1 U440 ( .A(G122), .B(G140), .ZN(n502) );
  INV_X1 U441 ( .A(KEYINPUT66), .ZN(n415) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n474) );
  INV_X1 U443 ( .A(KEYINPUT2), .ZN(n416) );
  NAND2_X1 U444 ( .A1(n414), .A2(n413), .ZN(n392) );
  INV_X1 U445 ( .A(n771), .ZN(n414) );
  XNOR2_X1 U446 ( .A(n419), .B(n418), .ZN(n437) );
  INV_X1 U447 ( .A(KEYINPUT25), .ZN(n418) );
  NAND2_X1 U448 ( .A1(n440), .A2(G217), .ZN(n419) );
  XNOR2_X1 U449 ( .A(n428), .B(n421), .ZN(n429) );
  XOR2_X1 U450 ( .A(G128), .B(G110), .Z(n421) );
  XNOR2_X1 U451 ( .A(G119), .B(G137), .ZN(n426) );
  XNOR2_X1 U452 ( .A(n491), .B(n360), .ZN(n649) );
  XNOR2_X1 U453 ( .A(n758), .B(n483), .ZN(n360) );
  NAND2_X1 U454 ( .A1(n600), .A2(n356), .ZN(n576) );
  NOR2_X1 U455 ( .A1(n541), .A2(n687), .ZN(n368) );
  OR2_X1 U456 ( .A1(n629), .A2(n687), .ZN(n473) );
  XNOR2_X1 U457 ( .A(n367), .B(n365), .ZN(n523) );
  NAND2_X1 U458 ( .A1(n521), .A2(G217), .ZN(n365) );
  AND2_X1 U459 ( .A1(n652), .A2(G953), .ZN(n755) );
  NAND2_X1 U460 ( .A1(n375), .A2(n374), .ZN(n373) );
  AND2_X1 U461 ( .A1(n554), .A2(n553), .ZN(n736) );
  AND2_X1 U462 ( .A1(n567), .A2(n529), .ZN(n738) );
  XOR2_X1 U463 ( .A(n449), .B(KEYINPUT97), .Z(n352) );
  XOR2_X1 U464 ( .A(G475), .B(n512), .Z(n353) );
  XOR2_X1 U465 ( .A(n593), .B(KEYINPUT81), .Z(n354) );
  OR2_X1 U466 ( .A1(n643), .A2(n642), .ZN(n355) );
  AND2_X1 U467 ( .A1(n738), .A2(n368), .ZN(n356) );
  AND2_X1 U468 ( .A1(n700), .A2(n695), .ZN(n357) );
  AND2_X1 U469 ( .A1(n594), .A2(KEYINPUT34), .ZN(n358) );
  NAND2_X2 U470 ( .A1(n376), .A2(n373), .ZN(n681) );
  AND2_X1 U471 ( .A1(n415), .A2(n416), .ZN(n359) );
  NAND2_X1 U472 ( .A1(n361), .A2(n357), .ZN(n604) );
  INV_X1 U473 ( .A(n605), .ZN(n601) );
  NAND2_X1 U474 ( .A1(n696), .A2(n547), .ZN(n457) );
  XNOR2_X2 U475 ( .A(n444), .B(n443), .ZN(n696) );
  XNOR2_X1 U476 ( .A(n575), .B(n574), .ZN(n364) );
  NAND2_X1 U477 ( .A1(n364), .A2(n779), .ZN(n363) );
  NAND2_X1 U478 ( .A1(n392), .A2(n359), .ZN(n391) );
  INV_X1 U479 ( .A(n621), .ZN(n361) );
  XNOR2_X2 U480 ( .A(n591), .B(n590), .ZN(n627) );
  NAND2_X1 U481 ( .A1(n684), .A2(n388), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n362), .A2(n610), .ZN(n617) );
  NAND2_X1 U483 ( .A1(n608), .A2(n609), .ZN(n362) );
  INV_X1 U484 ( .A(n369), .ZN(n409) );
  NAND2_X1 U485 ( .A1(n369), .A2(n546), .ZN(n401) );
  NAND2_X1 U486 ( .A1(n411), .A2(n410), .ZN(n369) );
  AND2_X2 U487 ( .A1(n370), .A2(n355), .ZN(n645) );
  AND2_X1 U488 ( .A1(n370), .A2(KEYINPUT82), .ZN(n413) );
  NAND2_X1 U489 ( .A1(n370), .A2(n772), .ZN(n761) );
  XNOR2_X2 U490 ( .A(n396), .B(KEYINPUT45), .ZN(n370) );
  XNOR2_X2 U491 ( .A(n770), .B(n455), .ZN(n656) );
  XNOR2_X2 U492 ( .A(n467), .B(n352), .ZN(n770) );
  XNOR2_X2 U493 ( .A(n522), .B(KEYINPUT4), .ZN(n488) );
  INV_X1 U494 ( .A(n695), .ZN(n582) );
  NAND2_X1 U495 ( .A1(n372), .A2(n415), .ZN(n390) );
  NAND2_X1 U496 ( .A1(n682), .A2(n417), .ZN(n372) );
  INV_X1 U497 ( .A(n382), .ZN(n375) );
  NAND2_X1 U498 ( .A1(n382), .A2(n594), .ZN(n377) );
  INV_X1 U499 ( .A(n594), .ZN(n378) );
  NAND2_X1 U500 ( .A1(n381), .A2(KEYINPUT34), .ZN(n379) );
  NAND2_X1 U501 ( .A1(n381), .A2(n358), .ZN(n380) );
  INV_X1 U502 ( .A(n686), .ZN(n381) );
  NOR2_X1 U503 ( .A1(n384), .A2(n354), .ZN(n383) );
  NOR2_X1 U504 ( .A1(n630), .A2(n592), .ZN(n384) );
  NAND2_X1 U505 ( .A1(n686), .A2(n386), .ZN(n385) );
  AND2_X1 U506 ( .A1(n630), .A2(n592), .ZN(n386) );
  NAND2_X1 U507 ( .A1(n392), .A2(n416), .ZN(n684) );
  XNOR2_X1 U508 ( .A(n393), .B(KEYINPUT113), .ZN(n565) );
  XNOR2_X2 U509 ( .A(n395), .B(KEYINPUT10), .ZN(n769) );
  XNOR2_X2 U510 ( .A(G146), .B(G125), .ZN(n395) );
  NAND2_X1 U511 ( .A1(n645), .A2(n644), .ZN(n682) );
  XNOR2_X2 U512 ( .A(n461), .B(n460), .ZN(n482) );
  OR2_X1 U513 ( .A1(n656), .A2(n406), .ZN(n405) );
  INV_X1 U514 ( .A(n397), .ZN(n404) );
  NAND2_X1 U515 ( .A1(n401), .A2(n398), .ZN(n397) );
  OR2_X1 U516 ( .A1(n656), .A2(n399), .ZN(n398) );
  NAND2_X1 U517 ( .A1(n409), .A2(n405), .ZN(n547) );
  NAND2_X1 U518 ( .A1(n403), .A2(n409), .ZN(n402) );
  AND2_X1 U519 ( .A1(n405), .A2(KEYINPUT1), .ZN(n403) );
  NAND2_X1 U520 ( .A1(n656), .A2(G469), .ZN(n411) );
  INV_X1 U521 ( .A(n646), .ZN(n417) );
  BUF_X1 U522 ( .A(n686), .Z(n717) );
  XNOR2_X1 U523 ( .A(n769), .B(n425), .ZN(n430) );
  XOR2_X1 U524 ( .A(n498), .B(KEYINPUT75), .Z(n422) );
  AND2_X1 U525 ( .A1(n570), .A2(n735), .ZN(n423) );
  AND2_X1 U526 ( .A1(n571), .A2(n423), .ZN(n572) );
  XNOR2_X1 U527 ( .A(n484), .B(G146), .ZN(n486) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n574) );
  INV_X1 U529 ( .A(KEYINPUT7), .ZN(n516) );
  BUF_X1 U530 ( .A(n602), .Z(n695) );
  XNOR2_X1 U531 ( .A(n499), .B(n422), .ZN(n530) );
  XNOR2_X1 U532 ( .A(G134), .B(KEYINPUT118), .ZN(n528) );
  XNOR2_X1 U533 ( .A(n424), .B(G140), .ZN(n449) );
  INV_X1 U534 ( .A(n449), .ZN(n425) );
  XOR2_X1 U535 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U536 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U537 ( .A(n429), .B(n430), .ZN(n433) );
  NAND2_X1 U538 ( .A1(G234), .A2(n772), .ZN(n431) );
  NAND2_X1 U539 ( .A1(G221), .A2(n521), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n433), .B(n432), .ZN(n752) );
  NOR2_X1 U541 ( .A1(G902), .A2(n752), .ZN(n439) );
  XNOR2_X2 U542 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n434) );
  XNOR2_X2 U543 ( .A(n434), .B(n407), .ZN(n646) );
  XNOR2_X1 U544 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n435) );
  XOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT80), .Z(n436) );
  XNOR2_X1 U546 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X2 U547 ( .A(n439), .B(n438), .ZN(n700) );
  NAND2_X1 U548 ( .A1(G221), .A2(n440), .ZN(n442) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT21), .Z(n441) );
  XOR2_X1 U550 ( .A(n442), .B(n441), .Z(n699) );
  NOR2_X2 U551 ( .A1(n700), .A2(n699), .ZN(n444) );
  INV_X1 U552 ( .A(KEYINPUT71), .ZN(n443) );
  XNOR2_X2 U553 ( .A(n446), .B(n445), .ZN(n522) );
  XNOR2_X1 U554 ( .A(n447), .B(G137), .ZN(n448) );
  XNOR2_X1 U555 ( .A(n450), .B(G107), .ZN(n756) );
  INV_X1 U556 ( .A(KEYINPUT74), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n464), .B(n451), .ZN(n452) );
  XNOR2_X1 U558 ( .A(n756), .B(n452), .ZN(n483) );
  NAND2_X1 U559 ( .A1(n772), .A2(G227), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n453), .B(G146), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n483), .B(n454), .ZN(n455) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n456) );
  XOR2_X1 U563 ( .A(KEYINPUT73), .B(G119), .Z(n460) );
  NAND2_X1 U564 ( .A1(n506), .A2(G210), .ZN(n463) );
  XNOR2_X1 U565 ( .A(G146), .B(KEYINPUT5), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U568 ( .A(n482), .B(n466), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n468), .B(n467), .ZN(n674) );
  INV_X1 U570 ( .A(KEYINPUT76), .ZN(n469) );
  XNOR2_X1 U571 ( .A(n469), .B(G472), .ZN(n470) );
  NAND2_X1 U572 ( .A1(G214), .A2(n492), .ZN(n472) );
  XOR2_X1 U573 ( .A(KEYINPUT94), .B(n472), .Z(n687) );
  XNOR2_X1 U574 ( .A(n473), .B(KEYINPUT30), .ZN(n480) );
  XOR2_X1 U575 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n475) );
  XNOR2_X1 U576 ( .A(n475), .B(n474), .ZN(n477) );
  NAND2_X1 U577 ( .A1(G952), .A2(n477), .ZN(n714) );
  NOR2_X1 U578 ( .A1(G953), .A2(n714), .ZN(n587) );
  NAND2_X1 U579 ( .A1(n477), .A2(n476), .ZN(n584) );
  XNOR2_X1 U580 ( .A(KEYINPUT110), .B(n584), .ZN(n478) );
  NOR2_X1 U581 ( .A1(G900), .A2(n478), .ZN(n479) );
  NOR2_X1 U582 ( .A1(n587), .A2(n479), .ZN(n533) );
  NOR2_X1 U583 ( .A1(n480), .A2(n533), .ZN(n564) );
  NAND2_X1 U584 ( .A1(G224), .A2(n772), .ZN(n485) );
  XNOR2_X1 U585 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U586 ( .A(n487), .B(KEYINPUT17), .Z(n490) );
  INV_X1 U587 ( .A(n488), .ZN(n489) );
  XNOR2_X1 U588 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U589 ( .A1(n649), .A2(n646), .ZN(n494) );
  AND2_X1 U590 ( .A1(G210), .A2(n492), .ZN(n493) );
  INV_X1 U591 ( .A(n550), .ZN(n579) );
  INV_X1 U592 ( .A(KEYINPUT38), .ZN(n495) );
  XNOR2_X1 U593 ( .A(n579), .B(n495), .ZN(n688) );
  INV_X1 U594 ( .A(n688), .ZN(n496) );
  AND2_X1 U595 ( .A1(n564), .A2(n496), .ZN(n497) );
  NAND2_X1 U596 ( .A1(n565), .A2(n497), .ZN(n499) );
  XNOR2_X1 U597 ( .A(KEYINPUT39), .B(KEYINPUT88), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n501), .B(n500), .ZN(n505) );
  XOR2_X1 U599 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n503) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U601 ( .A(n505), .B(n504), .Z(n511) );
  NAND2_X1 U602 ( .A1(G214), .A2(n506), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U604 ( .A(n509), .B(n769), .ZN(n510) );
  XNOR2_X1 U605 ( .A(n511), .B(n510), .ZN(n666) );
  NOR2_X1 U606 ( .A1(G902), .A2(n666), .ZN(n512) );
  INV_X1 U607 ( .A(KEYINPUT13), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n353), .B(n513), .ZN(n567) );
  XNOR2_X1 U609 ( .A(KEYINPUT107), .B(G478), .ZN(n526) );
  XNOR2_X1 U610 ( .A(n515), .B(n514), .ZN(n519) );
  XOR2_X1 U611 ( .A(n520), .B(KEYINPUT9), .Z(n524) );
  XNOR2_X1 U612 ( .A(n524), .B(n523), .ZN(n748) );
  NOR2_X1 U613 ( .A1(G902), .A2(n748), .ZN(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n566) );
  INV_X1 U615 ( .A(n566), .ZN(n529) );
  NOR2_X1 U616 ( .A1(n567), .A2(n529), .ZN(n527) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT108), .ZN(n741) );
  AND2_X1 U618 ( .A1(n530), .A2(n741), .ZN(n640) );
  XOR2_X1 U619 ( .A(n528), .B(n640), .Z(G36) );
  NAND2_X1 U620 ( .A1(n530), .A2(n738), .ZN(n531) );
  NOR2_X1 U621 ( .A1(n687), .A2(n688), .ZN(n691) );
  NOR2_X1 U622 ( .A1(n566), .A2(n567), .ZN(n689) );
  NAND2_X1 U623 ( .A1(n691), .A2(n689), .ZN(n532) );
  XNOR2_X1 U624 ( .A(KEYINPUT41), .B(n532), .ZN(n716) );
  INV_X1 U625 ( .A(n699), .ZN(n596) );
  INV_X1 U626 ( .A(n700), .ZN(n622) );
  NAND2_X1 U627 ( .A1(n596), .A2(n534), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n535), .B(KEYINPUT28), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n716), .A2(n554), .ZN(n537) );
  XNOR2_X1 U630 ( .A(n537), .B(KEYINPUT42), .ZN(n781) );
  NAND2_X1 U631 ( .A1(n673), .A2(n781), .ZN(n540) );
  XNOR2_X1 U632 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n538), .B(KEYINPUT64), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n540), .B(n539), .ZN(n573) );
  INV_X1 U635 ( .A(n687), .ZN(n549) );
  INV_X1 U636 ( .A(KEYINPUT109), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n542), .B(KEYINPUT6), .ZN(n543) );
  XNOR2_X1 U638 ( .A(n629), .B(n543), .ZN(n600) );
  INV_X1 U639 ( .A(n600), .ZN(n544) );
  NOR2_X1 U640 ( .A1(n579), .A2(n576), .ZN(n545) );
  XOR2_X1 U641 ( .A(KEYINPUT36), .B(n545), .Z(n548) );
  INV_X1 U642 ( .A(KEYINPUT1), .ZN(n546) );
  NOR2_X1 U643 ( .A1(n548), .A2(n582), .ZN(n744) );
  INV_X1 U644 ( .A(n589), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n736), .A2(KEYINPUT78), .ZN(n555) );
  NAND2_X1 U646 ( .A1(n555), .A2(KEYINPUT47), .ZN(n558) );
  OR2_X1 U647 ( .A1(n741), .A2(n738), .ZN(n560) );
  INV_X1 U648 ( .A(n560), .ZN(n632) );
  NAND2_X1 U649 ( .A1(n632), .A2(KEYINPUT47), .ZN(n556) );
  XOR2_X1 U650 ( .A(n556), .B(KEYINPUT83), .Z(n557) );
  NAND2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U652 ( .A1(n744), .A2(n559), .ZN(n571) );
  AND2_X1 U653 ( .A1(n560), .A2(n736), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n561), .B(KEYINPUT78), .ZN(n563) );
  INV_X1 U655 ( .A(KEYINPUT47), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n563), .A2(n562), .ZN(n570) );
  AND2_X1 U657 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U658 ( .A1(n567), .A2(n566), .ZN(n593) );
  NOR2_X1 U659 ( .A1(n579), .A2(n593), .ZN(n568) );
  NAND2_X1 U660 ( .A1(n569), .A2(n568), .ZN(n735) );
  NAND2_X1 U661 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U662 ( .A(KEYINPUT111), .B(n576), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n577), .A2(n582), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n578), .B(KEYINPUT43), .ZN(n580) );
  NAND2_X1 U665 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U666 ( .A(n581), .B(KEYINPUT112), .ZN(n779) );
  NAND2_X1 U667 ( .A1(n625), .A2(n600), .ZN(n583) );
  NOR2_X1 U668 ( .A1(G898), .A2(n584), .ZN(n585) );
  XNOR2_X1 U669 ( .A(n585), .B(KEYINPUT96), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X2 U671 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U672 ( .A(KEYINPUT0), .ZN(n590) );
  INV_X1 U673 ( .A(n627), .ZN(n630) );
  INV_X1 U674 ( .A(KEYINPUT34), .ZN(n592) );
  XNOR2_X1 U675 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n594) );
  XNOR2_X1 U676 ( .A(n681), .B(KEYINPUT70), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT77), .B(n595), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n689), .A2(n596), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n601), .A2(n544), .ZN(n621) );
  INV_X1 U681 ( .A(KEYINPUT32), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n622), .A2(n605), .ZN(n606) );
  AND2_X1 U683 ( .A1(n629), .A2(n606), .ZN(n607) );
  AND2_X1 U684 ( .A1(n582), .A2(n607), .ZN(n731) );
  NOR2_X1 U685 ( .A1(n780), .A2(n731), .ZN(n608) );
  INV_X1 U686 ( .A(KEYINPUT44), .ZN(n610) );
  INV_X1 U687 ( .A(n681), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n618), .A2(KEYINPUT90), .ZN(n615) );
  INV_X1 U689 ( .A(n731), .ZN(n612) );
  AND2_X1 U690 ( .A1(KEYINPUT70), .A2(KEYINPUT44), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n780), .A2(n613), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n638) );
  NAND2_X1 U695 ( .A1(n618), .A2(KEYINPUT44), .ZN(n620) );
  INV_X1 U696 ( .A(KEYINPUT90), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n636) );
  XOR2_X1 U698 ( .A(KEYINPUT89), .B(n621), .Z(n624) );
  NAND2_X1 U699 ( .A1(n582), .A2(n622), .ZN(n623) );
  BUF_X1 U700 ( .A(n625), .Z(n626) );
  INV_X1 U701 ( .A(n629), .ZN(n702) );
  NAND2_X1 U702 ( .A1(n626), .A2(n702), .ZN(n706) );
  NOR2_X1 U703 ( .A1(n706), .A2(n627), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT31), .B(n628), .Z(n740) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  OR2_X1 U706 ( .A1(n740), .A2(n412), .ZN(n633) );
  AND2_X1 U707 ( .A1(n633), .A2(n560), .ZN(n634) );
  NOR2_X1 U708 ( .A1(n725), .A2(n634), .ZN(n635) );
  AND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n643) );
  INV_X1 U712 ( .A(n640), .ZN(n641) );
  NOR2_X1 U713 ( .A1(n641), .A2(KEYINPUT82), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n747), .A2(G210), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n647) );
  XOR2_X1 U716 ( .A(n647), .B(KEYINPUT55), .Z(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n651), .B(n650), .ZN(n653) );
  INV_X1 U719 ( .A(G952), .ZN(n652) );
  INV_X1 U720 ( .A(n755), .ZN(n677) );
  NAND2_X1 U721 ( .A1(n653), .A2(n677), .ZN(n655) );
  INV_X1 U722 ( .A(KEYINPUT56), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n747), .A2(G469), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT123), .B(KEYINPUT122), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n656), .B(n659), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n662), .A2(n677), .ZN(n664) );
  INV_X1 U731 ( .A(KEYINPUT124), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(G54) );
  NAND2_X1 U733 ( .A1(n747), .A2(G475), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT68), .B(KEYINPUT59), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n669), .A2(n677), .ZN(n671) );
  INV_X1 U738 ( .A(KEYINPUT60), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G60) );
  XOR2_X1 U740 ( .A(G131), .B(KEYINPUT127), .Z(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(G33) );
  NAND2_X1 U742 ( .A1(n747), .A2(G472), .ZN(n676) );
  XOR2_X1 U743 ( .A(n674), .B(KEYINPUT62), .Z(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n679) );
  XNOR2_X1 U747 ( .A(n680), .B(n679), .ZN(G57) );
  XNOR2_X1 U748 ( .A(n681), .B(G122), .ZN(G24) );
  BUF_X1 U749 ( .A(n682), .Z(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT84), .ZN(n722) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U754 ( .A1(n691), .A2(n560), .ZN(n692) );
  NAND2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n717), .A2(n694), .ZN(n711) );
  XOR2_X1 U757 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n698) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U759 ( .A(n698), .B(n697), .Z(n705) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(KEYINPUT49), .B(n701), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U763 ( .A1(n705), .A2(n704), .ZN(n707) );
  AND2_X1 U764 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U765 ( .A(KEYINPUT51), .B(n708), .ZN(n709) );
  NAND2_X1 U766 ( .A1(n716), .A2(n709), .ZN(n710) );
  NAND2_X1 U767 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U768 ( .A(KEYINPUT52), .B(n712), .Z(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n715), .B(KEYINPUT120), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U772 ( .A1(n718), .A2(n772), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U775 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n724), .B(n723), .ZN(G75) );
  XOR2_X1 U777 ( .A(n725), .B(G101), .Z(G3) );
  NAND2_X1 U778 ( .A1(n412), .A2(n738), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n726), .B(G104), .ZN(G6) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT27), .ZN(n730) );
  XOR2_X1 U781 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n728) );
  NAND2_X1 U782 ( .A1(n412), .A2(n741), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n730), .B(n729), .ZN(G9) );
  XNOR2_X1 U785 ( .A(n731), .B(G110), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n732), .B(KEYINPUT115), .ZN(G12) );
  XOR2_X1 U787 ( .A(G128), .B(KEYINPUT29), .Z(n734) );
  NAND2_X1 U788 ( .A1(n736), .A2(n741), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n734), .B(n733), .ZN(G30) );
  XNOR2_X1 U790 ( .A(G143), .B(n735), .ZN(G45) );
  NAND2_X1 U791 ( .A1(n736), .A2(n738), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n737), .B(G146), .ZN(G48) );
  NAND2_X1 U793 ( .A1(n740), .A2(n738), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n739), .B(G113), .ZN(G15) );
  NAND2_X1 U795 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(KEYINPUT116), .ZN(n743) );
  XNOR2_X1 U797 ( .A(G116), .B(n743), .ZN(G18) );
  XOR2_X1 U798 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n746) );
  XNOR2_X1 U799 ( .A(n744), .B(G125), .ZN(n745) );
  XNOR2_X1 U800 ( .A(n746), .B(n745), .ZN(G27) );
  NAND2_X1 U801 ( .A1(n751), .A2(G478), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U803 ( .A1(n755), .A2(n750), .ZN(G63) );
  NAND2_X1 U804 ( .A1(n751), .A2(G217), .ZN(n753) );
  XNOR2_X1 U805 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(G66) );
  XOR2_X1 U807 ( .A(G101), .B(n756), .Z(n757) );
  XNOR2_X1 U808 ( .A(n758), .B(n757), .ZN(n760) );
  NOR2_X1 U809 ( .A1(G898), .A2(n772), .ZN(n759) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n768) );
  XNOR2_X1 U811 ( .A(n761), .B(KEYINPUT126), .ZN(n766) );
  XOR2_X1 U812 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n763) );
  NAND2_X1 U813 ( .A1(G224), .A2(G953), .ZN(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(n764) );
  NAND2_X1 U815 ( .A1(n764), .A2(G898), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U817 ( .A(n768), .B(n767), .ZN(G69) );
  XNOR2_X1 U818 ( .A(n770), .B(n769), .ZN(n774) );
  XNOR2_X1 U819 ( .A(n771), .B(n774), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(n772), .ZN(n778) );
  XNOR2_X1 U821 ( .A(n774), .B(G227), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n776), .A2(G953), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n778), .A2(n777), .ZN(G72) );
  XNOR2_X1 U825 ( .A(G140), .B(n779), .ZN(G42) );
  XOR2_X1 U826 ( .A(n780), .B(G119), .Z(G21) );
  XNOR2_X1 U827 ( .A(G137), .B(n781), .ZN(G39) );
endmodule

