//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G50), .A2(G226), .ZN(new_n209));
  AND2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n215), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G77), .A2(G244), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n207), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(new_n203), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n207), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  NOR3_X1   g0034(.A1(new_n225), .A2(new_n229), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n217), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n211), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  OAI21_X1  g0052(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n227), .A2(G33), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n228), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n262), .B1(new_n246), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(new_n263), .B2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n246), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G223), .A2(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n271), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n281), .C1(G77), .C2(new_n274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n283), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n282), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT67), .B(G179), .Z(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n269), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n269), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n266), .B(KEYINPUT9), .C1(new_n246), .C2(new_n268), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(G200), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n297), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT70), .B(KEYINPUT10), .Z(new_n304));
  OR3_X1    g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n310), .A3(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n295), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n280), .A2(G238), .A3(new_n283), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n271), .A2(new_n213), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G226), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n212), .B2(G1698), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n317), .B2(new_n274), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n286), .B(new_n314), .C1(new_n318), .C2(new_n280), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n212), .A2(G1698), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G226), .B2(G1698), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n322), .A2(new_n325), .B1(new_n271), .B2(new_n213), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n281), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n286), .A4(new_n314), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G179), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT76), .B(KEYINPUT14), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n330), .A2(KEYINPUT75), .A3(G169), .A4(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n336));
  AOI221_X4 g0136(.A(new_n292), .B1(new_n335), .B2(new_n336), .C1(new_n320), .C2(new_n329), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n332), .B(new_n334), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n341));
  AOI22_X1  g0141(.A1(G68), .A2(new_n267), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n256), .A2(new_n246), .B1(new_n227), .B2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(G77), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n259), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n262), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n264), .A2(G77), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n257), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT15), .B(G87), .Z(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n259), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n356), .B2(new_n262), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n344), .B2(new_n268), .ZN(new_n358));
  INV_X1    g0158(.A(G244), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n281), .B1(new_n274), .B2(G107), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G238), .A2(G1698), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n212), .B2(G1698), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n325), .A2(new_n362), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n286), .B1(new_n288), .B2(new_n359), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n358), .B1(new_n367), .B2(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n290), .B1(new_n365), .B2(new_n366), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g0170(.A(new_n364), .B(KEYINPUT68), .Z(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n298), .ZN(new_n372));
  INV_X1    g0172(.A(new_n358), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n351), .B1(new_n376), .B2(KEYINPUT69), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n280), .A2(G232), .A3(new_n283), .ZN(new_n379));
  OR2_X1    g0179(.A1(G223), .A2(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n287), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n323), .C2(new_n324), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n286), .B(new_n379), .C1(new_n384), .C2(new_n280), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G190), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n385), .B(KEYINPUT79), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n374), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n257), .A2(new_n265), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n268), .B2(new_n257), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n272), .A2(new_n227), .A3(new_n273), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n273), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(KEYINPUT77), .A3(new_n393), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G68), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n211), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n202), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT78), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n255), .A2(G159), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT78), .B(G20), .C1(new_n401), .C2(new_n202), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n400), .B1(new_n394), .B2(new_n396), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n262), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n391), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n388), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT17), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n413), .A2(new_n262), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n390), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n280), .B1(new_n382), .B2(new_n383), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n285), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n379), .ZN(new_n423));
  INV_X1    g0223(.A(new_n379), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n421), .A2(new_n424), .A3(KEYINPUT79), .A4(new_n285), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n419), .B1(new_n427), .B2(new_n386), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n292), .B1(new_n423), .B2(new_n425), .ZN(new_n433));
  INV_X1    g0233(.A(new_n290), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n422), .A2(new_n434), .A3(new_n379), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n415), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n415), .A3(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n378), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n441), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(new_n431), .A3(KEYINPUT80), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n313), .B(new_n377), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n376), .A2(KEYINPUT69), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n330), .A2(G200), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n349), .B1(new_n331), .B2(G190), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT74), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n445), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(new_n275), .C1(new_n323), .C2(new_n324), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(G250), .A2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n323), .B2(new_n324), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT82), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n459), .C1(new_n323), .C2(new_n324), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n461), .A2(new_n463), .B1(G33), .B2(G283), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n280), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(G274), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n469), .B2(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n280), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(new_n214), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT83), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n461), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n456), .A3(new_n457), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n281), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g0279(.A(new_n473), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n481), .A3(new_n292), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n434), .A3(new_n480), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT7), .B1(new_n325), .B2(new_n227), .ZN(new_n484));
  INV_X1    g0284(.A(new_n396), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g0286(.A(KEYINPUT81), .B(G107), .Z(new_n487));
  OR2_X1    g0287(.A1(KEYINPUT6), .A2(G97), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT81), .B(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n489), .A3(new_n488), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(G20), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n255), .A2(G77), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n262), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n261), .A2(new_n228), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n264), .C1(G1), .C2(new_n271), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n265), .A2(new_n213), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n482), .A2(new_n483), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n298), .B1(new_n474), .B2(new_n481), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n465), .B2(new_n473), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n501), .A3(new_n502), .A4(new_n497), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT84), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n510));
  AOI211_X1 g0310(.A(KEYINPUT83), .B(new_n473), .C1(new_n477), .C2(new_n281), .ZN(new_n511));
  OAI21_X1  g0311(.A(G190), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n374), .B1(new_n478), .B2(new_n480), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n504), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n482), .A2(new_n483), .A3(new_n503), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT84), .B1(new_n505), .B2(new_n507), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n512), .A2(new_n514), .A3(new_n509), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT85), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n280), .B1(new_n325), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G264), .A2(G1698), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n214), .B2(G1698), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n325), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n471), .A2(G270), .A3(new_n280), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n470), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G179), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n261), .A2(new_n228), .B1(G20), .B2(new_n216), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n476), .B(new_n227), .C1(G33), .C2(new_n213), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(KEYINPUT90), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n533), .B(new_n534), .C1(KEYINPUT90), .C2(new_n536), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n265), .A2(G116), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n499), .B2(G116), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n530), .A2(G200), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n538), .A2(new_n539), .B1(KEYINPUT90), .B2(new_n536), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n544), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n550), .C1(new_n298), .C2(new_n530), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n530), .B(G169), .C1(new_n544), .C2(new_n549), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n546), .A2(KEYINPUT21), .A3(G169), .A4(new_n530), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n547), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n227), .B(G87), .C1(new_n323), .C2(new_n324), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT22), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n227), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT23), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n271), .A2(new_n216), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n227), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n558), .A2(KEYINPUT24), .A3(new_n560), .A4(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n262), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n500), .A2(G107), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n264), .A2(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT25), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n470), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n471), .A2(G264), .A3(new_n280), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n220), .A2(new_n275), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n214), .A2(G1698), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n323), .C2(new_n324), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n281), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT91), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n471), .A2(new_n581), .A3(G264), .A4(new_n280), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT92), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT92), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n574), .A2(new_n580), .A3(new_n585), .A4(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(G179), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n580), .A2(new_n470), .A3(new_n573), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(G169), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n571), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n587), .A2(G200), .B1(G190), .B2(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(G97), .A2(G107), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n227), .A2(new_n595), .B1(new_n596), .B2(new_n219), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n274), .A2(new_n227), .A3(G68), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n227), .A2(G33), .A3(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT89), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT89), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n262), .B1(new_n601), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n354), .A2(new_n264), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n500), .A2(new_n354), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n359), .A2(G1698), .ZN(new_n615));
  OAI221_X1 g0415(.A(new_n615), .B1(G238), .B2(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n281), .B1(new_n617), .B2(new_n561), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n220), .B1(new_n466), .B2(G1), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n263), .A2(new_n284), .A3(G45), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n280), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT86), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n280), .A2(new_n623), .A3(new_n619), .A4(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(new_n625), .A3(new_n434), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n618), .A2(new_n625), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n292), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n618), .A2(new_n625), .A3(KEYINPUT87), .A4(new_n434), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n614), .A2(new_n628), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n606), .A2(new_n608), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n602), .A3(new_n599), .A4(new_n600), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n611), .B1(new_n634), .B2(new_n262), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n618), .A2(new_n625), .A3(G190), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(G200), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n500), .A2(G87), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n556), .A2(new_n591), .A3(new_n594), .A4(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n453), .A2(new_n518), .A3(new_n523), .A4(new_n642), .ZN(G372));
  NAND3_X1  g0443(.A1(new_n614), .A2(new_n630), .A3(new_n626), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n519), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n504), .B2(new_n640), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT93), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n520), .A2(new_n521), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n645), .B1(new_n592), .B2(new_n593), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n554), .A2(new_n555), .A3(new_n547), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n590), .B1(new_n587), .B2(G179), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n592), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n504), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT93), .A4(new_n644), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n652), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n453), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT94), .ZN(new_n662));
  INV_X1    g0462(.A(new_n370), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n351), .B1(new_n663), .B2(new_n451), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n441), .B1(new_n664), .B2(new_n431), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n307), .A2(new_n312), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n295), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G369));
  NOR2_X1   g0468(.A1(new_n230), .A2(G20), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .A3(G1), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n670), .B2(G1), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n550), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT95), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n554), .A2(new_n555), .A3(new_n547), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n556), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n591), .B(new_n594), .C1(new_n592), .C2(new_n675), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n591), .B2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n675), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n591), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n678), .A2(new_n675), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT96), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n231), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR4_X1   g0495(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n226), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n660), .A2(new_n675), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT98), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n658), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n522), .A2(KEYINPUT98), .A3(new_n657), .A4(new_n654), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n504), .B2(new_n645), .ZN(new_n706));
  INV_X1    g0506(.A(new_n644), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n504), .A2(new_n640), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n647), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n704), .A2(new_n705), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n629), .B1(new_n584), .B2(new_n586), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n712), .B(new_n532), .C1(new_n510), .C2(new_n511), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n584), .A2(new_n586), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n528), .A2(new_n529), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n470), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n478), .A2(new_n480), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n434), .A3(new_n719), .A4(new_n629), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n474), .A2(new_n481), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n532), .A4(new_n712), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n723), .B2(new_n688), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT97), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n518), .A2(new_n523), .A3(new_n642), .A4(new_n675), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n726), .B(new_n727), .C1(new_n729), .C2(KEYINPUT97), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n702), .A2(new_n711), .B1(G330), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n699), .B1(new_n731), .B2(G1), .ZN(G364));
  AOI21_X1  g0532(.A(new_n228), .B1(G20), .B2(new_n292), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n434), .A2(new_n227), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n374), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT101), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n227), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n735), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n742), .A2(G68), .B1(G107), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n298), .A2(new_n374), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n734), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G50), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n734), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n734), .A2(KEYINPUT100), .A3(new_n751), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n298), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n531), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n756), .A2(G77), .B1(G97), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n746), .A2(new_n274), .A3(new_n750), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n743), .A2(new_n751), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n762), .A2(KEYINPUT32), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n747), .A2(new_n743), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n219), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT32), .B1(new_n762), .B2(new_n763), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n734), .A2(new_n757), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n211), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n761), .A2(new_n764), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n742), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n765), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G303), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n749), .A2(G326), .ZN(new_n775));
  INV_X1    g0575(.A(new_n762), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n274), .B1(new_n776), .B2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n777), .B1(new_n778), .B2(new_n744), .C1(new_n752), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n768), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(G322), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n772), .A2(new_n774), .A3(new_n775), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G294), .B2(new_n759), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n733), .B1(new_n770), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n263), .B1(new_n669), .B2(G45), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n694), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT102), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n682), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n248), .A2(G45), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n231), .A2(new_n274), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G45), .C2(new_n226), .ZN(new_n798));
  INV_X1    g0598(.A(G355), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n232), .A2(new_n274), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(G116), .B2(new_n232), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n792), .A2(new_n733), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n785), .A2(new_n794), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT103), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n684), .A2(new_n788), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G330), .B2(new_n681), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(G396));
  AOI21_X1  g0608(.A(new_n325), .B1(new_n776), .B2(G132), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n742), .A2(G150), .B1(G143), .B2(new_n781), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  INV_X1    g0611(.A(new_n756), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n748), .C1(new_n763), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT34), .Z(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G50), .B2(new_n773), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n759), .A2(G58), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n745), .A2(G68), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n809), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n742), .A2(G283), .B1(G303), .B2(new_n749), .ZN(new_n819));
  INV_X1    g0619(.A(G107), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n765), .A2(new_n820), .B1(new_n744), .B2(new_n219), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n325), .B1(new_n768), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(G97), .C2(new_n759), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n819), .B(new_n824), .C1(new_n779), .C2(new_n762), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n756), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n733), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n827), .A2(new_n788), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n733), .A2(new_n790), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n368), .A2(new_n369), .A3(new_n688), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n372), .A2(new_n375), .B1(new_n373), .B2(new_n675), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n370), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n828), .B1(G77), .B2(new_n830), .C1(new_n791), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n700), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n660), .A2(new_n675), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n730), .A2(G330), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n838), .B(new_n839), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n789), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n834), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT113), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n674), .B1(new_n433), .B2(new_n435), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n399), .A2(new_n407), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n410), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT106), .A3(new_n262), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT106), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n399), .B2(new_n407), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n498), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n847), .A2(new_n408), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n844), .B1(new_n851), .B2(new_n391), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n852), .B2(new_n416), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n415), .A2(new_n674), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n437), .A2(new_n428), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT107), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n859), .B(KEYINPUT37), .C1(new_n852), .C2(new_n416), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n854), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n673), .B1(new_n851), .B2(new_n391), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n443), .B2(new_n431), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT112), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n727), .A2(new_n729), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n688), .A2(new_n349), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n350), .A2(new_n451), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n349), .B(new_n688), .C1(new_n339), .C2(KEYINPUT74), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n833), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n867), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(KEYINPUT112), .B(new_n873), .C1(new_n727), .C2(new_n729), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n866), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n843), .B1(new_n877), .B2(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n868), .A2(new_n874), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n861), .A2(new_n863), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n873), .B1(new_n727), .B2(new_n729), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n867), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n855), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n417), .A2(KEYINPUT109), .A3(new_n430), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n441), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT109), .B1(new_n417), .B2(new_n430), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n856), .B(new_n857), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n884), .A2(KEYINPUT110), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT110), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n861), .A2(new_n863), .A3(new_n900), .A4(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n902), .A2(new_n889), .A3(new_n879), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n891), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n453), .A2(new_n868), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n453), .A2(new_n702), .A3(new_n711), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n667), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT111), .Z(new_n911));
  XNOR2_X1  g0711(.A(new_n908), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n443), .A2(new_n673), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n831), .B(KEYINPUT104), .Z(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n837), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n885), .A3(new_n872), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n902), .B2(KEYINPUT39), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n350), .A2(new_n688), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n913), .B(new_n919), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n912), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n263), .B2(new_n669), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n491), .A2(new_n493), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n227), .B(new_n228), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(G116), .C1(new_n929), .C2(new_n928), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n226), .A2(new_n344), .A3(new_n401), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n201), .A2(new_n400), .ZN(new_n934));
  OAI211_X1 g0734(.A(G1), .B(new_n230), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n503), .A2(new_n688), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n522), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n519), .A2(new_n688), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n692), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n687), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n940), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT44), .B1(new_n692), .B2(new_n940), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n945), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n684), .B(new_n686), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n691), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n731), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n731), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n694), .B(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n786), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT42), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n940), .A2(new_n959), .A3(new_n686), .A4(new_n691), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT114), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n940), .A2(new_n686), .A3(new_n691), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n504), .B1(new_n938), .B2(new_n591), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n675), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n635), .A2(new_n638), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n688), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n646), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n707), .A2(new_n967), .A3(new_n688), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n971), .B(KEYINPUT43), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT115), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT115), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n966), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT116), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n972), .A2(new_n975), .A3(KEYINPUT116), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n940), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n687), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n687), .A2(new_n983), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n985), .A3(new_n981), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n958), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n742), .A2(G159), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n756), .A2(new_n201), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n274), .B1(new_n765), .B2(new_n211), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G68), .B2(new_n759), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n745), .A2(G77), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n811), .B2(new_n762), .C1(new_n768), .C2(new_n254), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G143), .B2(new_n749), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n762), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n756), .A2(G283), .B1(G107), .B2(new_n759), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n524), .B2(new_n768), .C1(new_n779), .C2(new_n748), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G294), .C2(new_n742), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n745), .A2(G97), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n773), .A2(G116), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT46), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n995), .B1(new_n1004), .B2(new_n274), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n733), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n969), .A2(new_n793), .A3(new_n970), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n797), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n802), .B1(new_n232), .B2(new_n355), .C1(new_n243), .C2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n788), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n987), .A2(new_n1011), .ZN(G387));
  INV_X1    g0812(.A(new_n733), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n756), .A2(G303), .B1(G322), .B2(new_n749), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n779), .B2(new_n741), .C1(new_n996), .C2(new_n768), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT48), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n759), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n778), .B2(new_n1017), .C1(new_n822), .C2(new_n765), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n274), .B1(new_n776), .B2(G326), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n216), .C2(new_n744), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n274), .B1(new_n752), .B2(new_n400), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G159), .B2(new_n749), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n246), .B2(new_n768), .C1(new_n355), .C2(new_n1017), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n765), .A2(new_n344), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n741), .A2(new_n258), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n1001), .C1(new_n254), .C2(new_n762), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1013), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n793), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n788), .B1(new_n686), .B2(new_n1030), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n258), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT50), .B1(new_n258), .B2(G50), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n466), .A4(new_n696), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n400), .A2(new_n344), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n797), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT117), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n466), .B2(new_n240), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(G107), .B2(new_n232), .C1(new_n696), .C2(new_n800), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT118), .Z(new_n1040));
  INV_X1    g0840(.A(new_n802), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1029), .A2(new_n1031), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n787), .B2(new_n953), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n954), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n694), .B1(new_n953), .B2(new_n731), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  AOI21_X1  g0847(.A(new_n695), .B1(new_n951), .B2(new_n954), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n951), .B2(new_n954), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n983), .A2(new_n792), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT120), .Z(new_n1051));
  OAI22_X1  g0851(.A1(new_n779), .A2(new_n768), .B1(new_n748), .B2(new_n996), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT121), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n274), .B1(new_n776), .B2(G322), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n752), .B2(new_n822), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n765), .A2(new_n778), .B1(new_n744), .B2(new_n820), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n742), .C2(G303), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1054), .B(new_n1058), .C1(new_n216), .C2(new_n1017), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT51), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n254), .A2(new_n748), .B1(new_n768), .B2(new_n763), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n742), .A2(new_n201), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n776), .A2(G143), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1061), .A2(new_n1060), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n765), .A2(new_n400), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n274), .B1(new_n744), .B2(new_n219), .C1(new_n1017), .C2(new_n344), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n756), .C2(new_n257), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1013), .B1(new_n1059), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n797), .A2(new_n251), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1041), .B1(new_n231), .B2(G97), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n789), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1051), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n951), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n949), .A2(KEYINPUT119), .A3(new_n950), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n787), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1049), .A2(new_n1073), .A3(new_n1077), .ZN(G390));
  NAND3_X1  g0878(.A1(new_n453), .A2(G330), .A3(new_n868), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n909), .A2(new_n1079), .A3(new_n667), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n879), .A2(new_n683), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n835), .A2(new_n683), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n872), .B1(new_n730), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n918), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n868), .A2(new_n1082), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n871), .A3(new_n870), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n730), .A2(new_n872), .A3(new_n1082), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n710), .A2(new_n675), .A3(new_n833), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n914), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1080), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1085), .A2(KEYINPUT122), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1088), .A2(new_n914), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n922), .B1(new_n1094), .B2(new_n872), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n899), .A2(new_n901), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n898), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n918), .A2(new_n872), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n923), .ZN(new_n1100));
  AOI221_X4 g0900(.A(new_n1093), .B1(new_n1095), .B2(new_n1098), .C1(new_n921), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1081), .A2(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n921), .A2(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1091), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1104), .C1(new_n1092), .C2(new_n1087), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1090), .B(new_n1107), .C1(new_n1108), .C2(new_n1102), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n694), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n921), .A2(new_n790), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n773), .A2(G150), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n742), .A2(G137), .B1(G159), .B2(new_n759), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n812), .B2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT123), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n776), .A2(G125), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G128), .A2(new_n749), .B1(new_n781), .B2(G132), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1118), .A2(new_n274), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1113), .B(new_n1121), .C1(new_n201), .C2(new_n745), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n756), .A2(G97), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n742), .A2(G107), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n781), .A2(G116), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n325), .B1(new_n748), .B2(new_n778), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n817), .B1(new_n822), .B2(new_n762), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(KEYINPUT124), .B1(new_n344), .B2(new_n1017), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .A4(new_n766), .ZN(new_n1130));
  AND4_X1   g0930(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n733), .B1(new_n1122), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1111), .A2(new_n788), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n258), .B2(new_n829), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n787), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1110), .A2(new_n1136), .ZN(G378));
  AND3_X1   g0937(.A1(new_n888), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT113), .B1(new_n888), .B2(new_n889), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n904), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT126), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n313), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n313), .A2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n269), .A2(new_n674), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1147), .A2(new_n1150), .A3(new_n1148), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1140), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n891), .A2(G330), .A3(new_n1154), .A4(new_n904), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1156), .A2(new_n925), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n925), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n787), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n325), .B1(new_n778), .B2(new_n762), .C1(new_n748), .C2(new_n216), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1025), .B1(G68), .B2(new_n759), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n211), .B2(new_n744), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n279), .B1(new_n768), .B2(new_n820), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n213), .B2(new_n741), .C1(new_n355), .C2(new_n752), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT58), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n246), .B1(new_n323), .B2(G41), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1017), .A2(new_n254), .B1(new_n765), .B2(new_n1116), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1170), .A2(new_n748), .B1(new_n752), .B2(new_n811), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n742), .C2(G132), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n768), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n1174), .B2(KEYINPUT59), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G33), .B1(new_n776), .B2(G124), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n763), .C2(new_n744), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1167), .B(new_n1168), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT125), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n789), .B1(new_n1180), .B2(new_n733), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n201), .B2(new_n830), .C1(new_n1154), .C2(new_n791), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1160), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n924), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT127), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1156), .A2(new_n1157), .A3(new_n925), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1159), .A2(KEYINPUT127), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1080), .B1(new_n1135), .B2(new_n1090), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1191), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n694), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1184), .B1(new_n1194), .B2(new_n1196), .ZN(G375));
  AOI21_X1  g0997(.A(new_n786), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n870), .A2(new_n790), .A3(new_n871), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n274), .B1(new_n752), .B2(new_n254), .C1(new_n811), .C2(new_n768), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n742), .B2(new_n1115), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1017), .A2(new_n246), .B1(new_n211), .B2(new_n744), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n749), .B2(G132), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n1173), .B2(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n812), .A2(new_n820), .B1(new_n822), .B2(new_n748), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n992), .B1(new_n213), .B2(new_n765), .C1(new_n1017), .C2(new_n355), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n325), .B1(new_n768), .B2(new_n778), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n216), .B2(new_n741), .C1(new_n524), .C2(new_n762), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1013), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n789), .B(new_n1211), .C1(new_n400), .C2(new_n829), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1198), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1080), .A2(new_n1084), .A3(new_n1089), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n956), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1213), .B1(new_n1215), .B2(new_n1090), .ZN(G381));
  INV_X1    g1016(.A(new_n1080), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1109), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n695), .B1(new_n1219), .B2(new_n1192), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1183), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1224), .A2(G384), .A3(G381), .ZN(new_n1225));
  INV_X1    g1025(.A(G390), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n987), .A3(new_n1011), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(G396), .A3(G393), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(G407));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1224), .ZN(G409));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1189), .A2(new_n787), .A3(new_n1190), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1195), .A2(new_n956), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1223), .A4(new_n1182), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n695), .B1(new_n1214), .B2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n1091), .C1(new_n1238), .C2(new_n1214), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1213), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n841), .A3(new_n834), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G384), .A2(new_n1240), .A3(new_n1213), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1232), .A2(G2897), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1237), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT63), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1232), .B1(G375), .B2(G378), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1244), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1236), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(G396), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1227), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1226), .B1(new_n987), .B2(new_n1011), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1227), .A3(new_n1254), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1237), .A2(new_n1244), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(KEYINPUT63), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1252), .A2(new_n1253), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1249), .A2(new_n1265), .A3(new_n1250), .A4(new_n1236), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT62), .B1(new_n1237), .B2(new_n1244), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1253), .A4(new_n1247), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1261), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(G405));
  NAND2_X1  g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1224), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(new_n1224), .A3(new_n1271), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1250), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1250), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G402));
endmodule


