//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  INV_X1    g000(.A(G127gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G134gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(G134gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G113gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(new_n208), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n208), .A2(G113gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n204), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n203), .A2(new_n205), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n207), .A2(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n219), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT27), .B(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n226), .A2(KEYINPUT28), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT28), .B1(new_n226), .B2(new_n227), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n233), .B2(new_n217), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n225), .A2(new_n235), .B1(new_n236), .B2(G190gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n225), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT25), .B1(new_n245), .B2(KEYINPUT65), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT23), .B1(new_n222), .B2(new_n223), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n218), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n248), .A3(new_n231), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n216), .B(new_n230), .C1(new_n242), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n230), .B1(new_n242), .B2(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n214), .A2(new_n215), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n209), .B1(new_n258), .B2(G120gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n255), .B1(new_n259), .B2(new_n206), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT64), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n241), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n249), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n216), .A4(new_n230), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n253), .A2(new_n261), .A3(new_n264), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT34), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n269), .B2(KEYINPUT71), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT32), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n261), .A3(new_n268), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n263), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n276), .B2(new_n263), .ZN(new_n280));
  XOR2_X1   g079(.A(G15gat), .B(G43gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT69), .ZN(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n277), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n278), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n287), .B2(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n277), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n274), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n277), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n263), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n278), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n284), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT34), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n271), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n299), .A3(new_n290), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n274), .C1(new_n286), .C2(new_n291), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT31), .B(G50gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G204gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G197gat), .ZN(new_n310));
  INV_X1    g109(.A(G197gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G204gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n313), .B(new_n314), .C1(new_n318), .C2(KEYINPUT22), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n314), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n310), .A2(new_n312), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n326));
  OAI21_X1  g125(.A(G218gat), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(KEYINPUT82), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n313), .B1(new_n318), .B2(KEYINPUT22), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n322), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n321), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT3), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  AND2_X1   g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(KEYINPUT77), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n339), .A2(new_n344), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n345), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n338), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT83), .B1(new_n335), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n345), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n346), .ZN(new_n361));
  INV_X1    g160(.A(new_n352), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n334), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n314), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G218gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n315), .A2(G211gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n331), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT74), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n375), .A2(KEYINPUT74), .B1(new_n367), .B2(new_n371), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n331), .A2(new_n373), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT76), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n319), .B(new_n365), .C1(new_n378), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n359), .A2(new_n363), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n319), .A2(new_n320), .B1(new_n331), .B2(new_n322), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n385), .B2(new_n330), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n384), .C1(new_n386), .C2(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n356), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G228gat), .A2(G233gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n377), .B1(new_n374), .B2(new_n376), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n379), .A2(KEYINPUT76), .A3(new_n380), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n391), .A2(new_n392), .B1(new_n329), .B2(new_n324), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n389), .B1(new_n393), .B2(new_n365), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n319), .B1(new_n378), .B2(new_n381), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n395), .B2(new_n334), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n396), .B2(new_n355), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n308), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n390), .A2(new_n397), .A3(new_n398), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n398), .B1(new_n390), .B2(new_n397), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT85), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  INV_X1    g205(.A(new_n389), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n384), .B1(new_n386), .B2(KEYINPUT3), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(KEYINPUT83), .B1(new_n393), .B2(new_n365), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n409), .B2(new_n387), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n382), .A2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n360), .B1(new_n393), .B2(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n384), .ZN(new_n413));
  OAI21_X1  g212(.A(G22gat), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n414), .B2(new_n399), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n402), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n254), .A2(new_n334), .B1(G226gat), .B2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n254), .A2(G226gat), .A3(G233gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n395), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n254), .A2(G226gat), .A3(G233gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n393), .B1(new_n421), .B2(new_n417), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n420), .A2(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT30), .A4(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT79), .B1(new_n384), .B2(new_n260), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n216), .A2(new_n355), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n384), .A2(new_n260), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT4), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT78), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(KEYINPUT3), .C1(new_n350), .C2(new_n354), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n364), .A3(new_n260), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT80), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n442), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n444), .A2(new_n364), .A3(new_n260), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT78), .B1(new_n355), .B2(new_n360), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n438), .A4(new_n440), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n216), .A2(new_n355), .A3(KEYINPUT81), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT81), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n384), .B2(new_n260), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n434), .B(new_n437), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n455), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n448), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n439), .A2(KEYINPUT4), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n434), .A2(new_n437), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT4), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n455), .A3(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G1gat), .B(G29gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT0), .ZN(new_n468));
  XNOR2_X1  g267(.A(G57gat), .B(G85gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(new_n470), .A3(new_n465), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n433), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT85), .B1(new_n403), .B2(new_n404), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n414), .A2(new_n406), .A3(new_n399), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n401), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n304), .A2(new_n416), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  INV_X1    g281(.A(new_n416), .ZN(new_n483));
  INV_X1    g282(.A(new_n480), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n292), .A2(new_n300), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(new_n477), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n482), .A2(KEYINPUT90), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n481), .A2(new_n490), .A3(KEYINPUT35), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n416), .A2(KEYINPUT86), .A3(new_n480), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT86), .B1(new_n416), .B2(new_n480), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n476), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n492), .A2(new_n493), .B1(new_n495), .B2(new_n433), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n450), .A2(new_n451), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n442), .B1(new_n464), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT39), .B1(new_n459), .B2(new_n449), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT39), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n470), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n500), .A2(KEYINPUT40), .A3(new_n470), .A4(new_n502), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n433), .A4(new_n472), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n416), .A2(new_n480), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n420), .B2(new_n422), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n510), .A2(new_n511), .A3(new_n425), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT88), .B1(new_n429), .B2(KEYINPUT37), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n420), .A2(new_n422), .A3(new_n514), .A4(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n510), .B2(new_n425), .ZN(new_n517));
  AND4_X1   g316(.A1(KEYINPUT38), .A2(new_n512), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n422), .A2(KEYINPUT87), .A3(new_n395), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n420), .A2(KEYINPUT87), .A3(new_n422), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n425), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT38), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n495), .B(new_n426), .C1(new_n518), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n486), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n304), .A2(KEYINPUT36), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n508), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n489), .A2(new_n491), .B1(new_n496), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G50gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT15), .B1(new_n530), .B2(G43gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(G43gat), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT14), .ZN(new_n534));
  INV_X1    g333(.A(G29gat), .ZN(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n532), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT92), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT93), .B(G43gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n530), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT94), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n530), .A2(G43gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n541), .A2(G50gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT15), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT95), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n537), .B(KEYINPUT96), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n551), .A2(new_n532), .A3(new_n534), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(KEYINPUT95), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n540), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT17), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT16), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(G1gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(G1gat), .B2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(G8gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n550), .A2(new_n552), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n539), .B1(new_n564), .B2(new_n554), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n556), .A2(new_n563), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n569), .A4(new_n570), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n556), .B(new_n563), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n569), .B(KEYINPUT13), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G169gat), .B(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT12), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n573), .A2(new_n574), .A3(new_n577), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n590), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n598), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n590), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n557), .A2(new_n567), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT103), .ZN(new_n605));
  INV_X1    g404(.A(new_n602), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n565), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n603), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n603), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G134gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n348), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n610), .B2(KEYINPUT104), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n611), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G71gat), .ZN(new_n618));
  INV_X1    g417(.A(G78gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G57gat), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n625), .A2(G64gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(G64gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT9), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(KEYINPUT99), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n624), .B2(new_n629), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT97), .B1(new_n618), .B2(new_n619), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n621), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n630), .A2(new_n631), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n563), .B1(new_n636), .B2(new_n637), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT101), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n644), .A3(new_n645), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n649), .A2(new_n655), .A3(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n636), .A2(new_n602), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  INV_X1    g463(.A(new_n601), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n636), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n636), .A2(new_n602), .A3(new_n664), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n663), .B1(new_n665), .B2(new_n636), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  OR2_X1    g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n662), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n617), .A2(new_n660), .A3(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n529), .A2(new_n589), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n495), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(G1gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1324gat));
  AND2_X1   g484(.A1(new_n682), .A2(new_n433), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n689), .B(new_n690), .C1(new_n562), .C2(new_n686), .ZN(G1325gat));
  AND2_X1   g490(.A1(new_n526), .A2(new_n527), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n682), .A2(G15gat), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n682), .A2(new_n525), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n492), .A2(new_n493), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NOR2_X1   g503(.A1(new_n529), .A2(new_n589), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n659), .A2(new_n680), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n617), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT107), .Z(new_n708));
  AND2_X1   g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n535), .A3(new_n495), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n706), .A2(new_n589), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n482), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n485), .A2(new_n488), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n491), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n528), .A2(new_n496), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n713), .B1(new_n718), .B2(new_n616), .ZN(new_n719));
  AOI211_X1 g518(.A(KEYINPUT44), .B(new_n617), .C1(new_n716), .C2(new_n717), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n712), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n494), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n711), .A2(new_n722), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n709), .A2(new_n536), .A3(new_n433), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT46), .Z(new_n725));
  INV_X1    g524(.A(new_n433), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1329gat));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n729), .A2(KEYINPUT109), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(KEYINPUT109), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n486), .A2(new_n542), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n705), .A2(new_n708), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT108), .ZN(new_n734));
  INV_X1    g533(.A(new_n712), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n529), .B2(new_n617), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n617), .B1(new_n716), .B2(new_n717), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n713), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n541), .B1(new_n739), .B2(new_n692), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n730), .B(new_n731), .C1(new_n734), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n733), .B(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n692), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n542), .B1(new_n721), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n743), .A2(new_n745), .A3(KEYINPUT109), .A4(new_n729), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n741), .A2(new_n746), .ZN(G1330gat));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n530), .B1(new_n739), .B2(new_n701), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n705), .A2(new_n530), .A3(new_n708), .A4(new_n701), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n748), .ZN(new_n753));
  OAI21_X1  g552(.A(G50gat), .B1(new_n721), .B2(new_n485), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(G1331gat));
  NOR4_X1   g557(.A1(new_n616), .A2(new_n659), .A3(new_n588), .A4(new_n680), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n718), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n494), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n625), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n726), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n760), .B2(new_n744), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n525), .A2(new_n618), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g570(.A1(new_n760), .A2(new_n700), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n619), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n589), .A2(new_n659), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n680), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n719), .B2(new_n720), .ZN(new_n777));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777), .B2(new_n494), .ZN(new_n778));
  INV_X1    g577(.A(new_n775), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n737), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n737), .A2(new_n779), .A3(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n495), .A2(new_n594), .A3(new_n679), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(G1336gat));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n680), .A2(new_n726), .A3(G92gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT112), .B2(new_n787), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n679), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n736), .B2(new_n738), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n595), .B1(new_n792), .B2(new_n433), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n788), .B(KEYINPUT113), .Z(new_n795));
  AOI22_X1  g594(.A1(new_n793), .A2(new_n794), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n790), .A2(new_n793), .B1(new_n796), .B2(new_n787), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n777), .B2(new_n744), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n680), .A2(G99gat), .A3(new_n486), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n784), .B2(new_n799), .ZN(G1338gat));
  NOR3_X1   g599(.A1(new_n485), .A2(G106gat), .A3(new_n680), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n780), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n485), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n792), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n701), .B(new_n776), .C1(new_n719), .C2(new_n720), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n804), .B1(new_n811), .B2(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n806), .B1(new_n792), .B2(new_n701), .ZN(new_n814));
  INV_X1    g613(.A(new_n801), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n781), .B2(new_n782), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n777), .B2(new_n485), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n804), .A3(new_n803), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n681), .A2(new_n588), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n666), .A2(new_n662), .A3(new_n667), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n676), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n827));
  AOI21_X1  g626(.A(new_n673), .B1(new_n668), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n678), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n828), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n588), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n575), .A2(new_n576), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n583), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n587), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n679), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n616), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n616), .A2(new_n839), .A3(new_n833), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n659), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n701), .A2(new_n486), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n494), .A2(new_n433), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n589), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n494), .B1(new_n824), .B2(new_n844), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n485), .A2(new_n304), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n433), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n258), .A3(new_n588), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n850), .A2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n208), .A3(new_n679), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n845), .A2(new_n679), .A3(new_n848), .A4(new_n846), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(G120gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(G120gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n849), .B2(new_n659), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n202), .A3(new_n660), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1342gat));
  OR3_X1    g666(.A1(new_n854), .A2(G134gat), .A3(new_n617), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n849), .B2(new_n617), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n744), .A2(new_n807), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n433), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n340), .B1(new_n875), .B2(new_n589), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n744), .A2(new_n848), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n485), .B1(new_n824), .B2(new_n844), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n832), .A2(new_n831), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT118), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n832), .A2(new_n883), .A3(new_n831), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n830), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n885), .A2(new_n588), .B1(new_n839), .B2(new_n679), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n886), .B2(new_n616), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n842), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n616), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n659), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n700), .B1(new_n890), .B2(new_n824), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n589), .A2(new_n340), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n876), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(new_n875), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n341), .A3(new_n679), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n842), .B1(new_n886), .B2(new_n616), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n660), .B1(new_n901), .B2(KEYINPUT121), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n823), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n700), .A2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n877), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n878), .A2(new_n879), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n907), .A2(new_n679), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n892), .A2(new_n680), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n900), .A2(G148gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n899), .B1(new_n911), .B2(new_n914), .ZN(G1345gat));
  OAI211_X1 g714(.A(new_n660), .B(new_n880), .C1(new_n891), .C2(new_n879), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G155gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n347), .A3(new_n660), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n892), .B2(new_n617), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n348), .A3(new_n616), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1347gat));
  AOI21_X1  g725(.A(new_n495), .B1(new_n824), .B2(new_n844), .ZN(new_n927));
  AND4_X1   g726(.A1(new_n433), .A2(new_n927), .A3(new_n485), .A4(new_n304), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n222), .A3(new_n588), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n494), .A2(new_n433), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n847), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n588), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT124), .B1(new_n934), .B2(G169gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n932), .B2(new_n680), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n928), .A2(new_n223), .A3(new_n679), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT125), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n932), .B2(new_n659), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n226), .A3(new_n660), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n227), .A3(new_n616), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n933), .A2(new_n616), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT61), .B(new_n227), .C1(new_n933), .C2(new_n616), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NAND2_X1  g750(.A1(new_n744), .A2(new_n931), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n909), .B(new_n953), .C1(new_n904), .C2(new_n906), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(new_n311), .A3(new_n589), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n873), .A2(new_n726), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n927), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n588), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n955), .A2(new_n959), .ZN(G1352gat));
  XNOR2_X1  g759(.A(KEYINPUT126), .B(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n907), .A2(new_n679), .A3(new_n909), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n952), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n957), .A2(new_n680), .A3(new_n961), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n368), .B1(KEYINPUT127), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n968), .B1(new_n954), .B2(new_n659), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT63), .ZN(new_n971));
  OAI221_X1 g770(.A(new_n968), .B1(KEYINPUT127), .B2(new_n967), .C1(new_n954), .C2(new_n659), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n958), .A2(new_n316), .A3(new_n317), .A4(new_n660), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n954), .B2(new_n617), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n315), .A3(new_n616), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


