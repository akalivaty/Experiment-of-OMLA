//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1148, new_n1149, new_n1150, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  AOI21_X1  g0049(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n250), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(new_n252), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n253), .B1(new_n255), .B2(G238), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n259), .B2(new_n231), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n260), .B1(G226), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n256), .B1(new_n267), .B2(new_n254), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G169), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT14), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT14), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n270), .A2(KEYINPUT14), .B1(new_n276), .B2(new_n269), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT66), .Z(new_n283));
  INV_X1    g0083(.A(new_n215), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n208), .B2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n206), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n244), .A2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n207), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n207), .A2(new_n262), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n290), .B1(new_n291), .B2(new_n219), .C1(new_n202), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n286), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n281), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(KEYINPUT12), .A3(new_n290), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n283), .A2(new_n244), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(KEYINPUT12), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n279), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n269), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n269), .A2(G200), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT8), .B(G58), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n309), .A2(new_n291), .B1(new_n310), .B2(new_n292), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G20), .B2(new_n203), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(new_n285), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n285), .A2(new_n282), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n288), .A2(G50), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n314), .A2(new_n315), .B1(G50), .B2(new_n282), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(KEYINPUT9), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT67), .ZN(new_n319));
  INV_X1    g0119(.A(new_n259), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G223), .B1(G77), .B2(new_n265), .ZN(new_n321));
  INV_X1    g0121(.A(G222), .ZN(new_n322));
  INV_X1    g0122(.A(new_n266), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n250), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n253), .B1(new_n255), .B2(G226), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G200), .B1(KEYINPUT9), .B2(new_n317), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n319), .B(new_n328), .C1(new_n304), .C2(new_n327), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT10), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n327), .A2(G179), .ZN(new_n331));
  INV_X1    g0131(.A(new_n317), .ZN(new_n332));
  INV_X1    g0132(.A(new_n327), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(G169), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n287), .A2(G77), .A3(new_n288), .ZN(new_n336));
  INV_X1    g0136(.A(new_n309), .ZN(new_n337));
  INV_X1    g0137(.A(new_n292), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(G20), .B2(G77), .ZN(new_n339));
  XOR2_X1   g0139(.A(KEYINPUT15), .B(G87), .Z(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n291), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n286), .B1(new_n283), .B2(new_n219), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n255), .A2(G244), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n320), .A2(G238), .B1(G107), .B2(new_n265), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n231), .B2(new_n323), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n253), .B(new_n345), .C1(new_n347), .C2(new_n250), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(G200), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n276), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n344), .C1(G169), .C2(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n308), .A2(new_n335), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n337), .A2(new_n288), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n314), .A2(new_n356), .B1(new_n282), .B2(new_n337), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n244), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n292), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT72), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n262), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT69), .A2(G33), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n261), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT70), .B1(new_n368), .B2(new_n264), .ZN(new_n369));
  AND2_X1   g0169(.A1(KEYINPUT69), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(KEYINPUT69), .A2(G33), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT3), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  INV_X1    g0173(.A(new_n264), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n207), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n374), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT71), .A3(G68), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n376), .B2(new_n377), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n244), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n364), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n366), .A2(new_n367), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n391), .A2(new_n380), .A3(new_n263), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n265), .B2(new_n207), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT73), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT73), .B(G68), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n363), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n285), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n357), .B1(new_n389), .B2(new_n400), .ZN(new_n401));
  MUX2_X1   g0201(.A(G223), .B(G226), .S(G1698), .Z(new_n402));
  AOI22_X1  g0202(.A1(new_n379), .A2(new_n402), .B1(G33), .B2(G87), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(new_n254), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n253), .B1(new_n255), .B2(G232), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G169), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT74), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n276), .A3(new_n405), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT18), .B1(new_n401), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n401), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n413), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n406), .A2(new_n304), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G200), .B2(new_n406), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n401), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n415), .A2(new_n418), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n355), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n207), .A2(G107), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT23), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n390), .A2(G116), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(G20), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G87), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n431), .A2(KEYINPUT22), .A3(G20), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n258), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g0233(.A(new_n433), .B(KEYINPUT80), .Z(new_n434));
  NAND3_X1  g0234(.A1(new_n379), .A2(new_n207), .A3(G87), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT22), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n430), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT24), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n285), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT25), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g0241(.A(new_n282), .ZN(new_n442));
  AOI21_X1  g0242(.A(G107), .B1(new_n440), .B2(KEYINPUT81), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n282), .A2(KEYINPUT81), .A3(new_n440), .A4(G107), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n285), .B(new_n282), .C1(G1), .C2(new_n262), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n444), .A2(new_n445), .B1(new_n446), .B2(new_n221), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n250), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G264), .ZN(new_n453));
  MUX2_X1   g0253(.A(G250), .B(G257), .S(G1698), .Z(new_n454));
  AOI22_X1  g0254(.A1(new_n379), .A2(new_n454), .B1(G294), .B2(new_n390), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n455), .B2(new_n254), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n250), .A2(new_n251), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n450), .A3(new_n451), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n456), .B(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n458), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(new_n276), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n448), .B1(KEYINPUT83), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n464), .A2(KEYINPUT83), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n221), .A3(KEYINPUT6), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(KEYINPUT6), .B2(new_n468), .ZN(new_n470));
  XOR2_X1   g0270(.A(KEYINPUT75), .B(G107), .Z(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(G20), .B1(G77), .B2(new_n338), .ZN(new_n473));
  OAI21_X1  g0273(.A(G107), .B1(new_n392), .B2(new_n393), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n285), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n442), .A2(new_n468), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n446), .B2(new_n468), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n459), .B1(G257), .B2(new_n452), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n320), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n368), .A2(new_n264), .ZN(new_n482));
  INV_X1    g0282(.A(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G244), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n479), .B1(new_n487), .B2(new_n254), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n276), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(G169), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n478), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n478), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(KEYINPUT76), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT76), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n488), .A2(new_n304), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(G200), .B2(new_n488), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n457), .A2(new_n450), .ZN(new_n501));
  OAI21_X1  g0301(.A(G250), .B1(new_n449), .B2(G1), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n250), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT77), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n220), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G238), .B2(G1698), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n429), .B1(new_n482), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n254), .B1(new_n507), .B2(KEYINPUT78), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(KEYINPUT78), .B2(new_n507), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n276), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n504), .A2(new_n509), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n407), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n379), .A2(new_n207), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n207), .B1(new_n257), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n431), .A2(new_n468), .A3(new_n221), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n516), .A2(new_n517), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n285), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n283), .B2(new_n341), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n341), .B2(new_n446), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n511), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n512), .A2(G200), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n446), .A2(new_n431), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n526), .C1(new_n304), .C2(new_n512), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n500), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n463), .A2(new_n350), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G190), .B2(new_n460), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n448), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n207), .C1(G33), .C2(new_n468), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT79), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n286), .C1(new_n207), .C2(G116), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT20), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G116), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n206), .B2(G33), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n287), .A2(new_n542), .B1(new_n541), .B2(new_n283), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n459), .B1(G270), .B2(new_n452), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n222), .A2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G257), .B2(G1698), .ZN(new_n547));
  INV_X1    g0347(.A(G303), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n482), .A2(new_n547), .B1(new_n548), .B2(new_n258), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n250), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G169), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n534), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n540), .A2(new_n543), .ZN(new_n554));
  INV_X1    g0354(.A(new_n551), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(G179), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n554), .A2(KEYINPUT21), .A3(G169), .A4(new_n551), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n554), .B1(G200), .B2(new_n551), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n304), .B2(new_n551), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR4_X1   g0361(.A1(new_n467), .A2(new_n529), .A3(new_n533), .A4(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n426), .A2(new_n562), .ZN(G372));
  INV_X1    g0363(.A(new_n330), .ZN(new_n564));
  INV_X1    g0364(.A(new_n307), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n303), .B1(new_n565), .B2(new_n353), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n423), .A2(new_n424), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n418), .A2(new_n415), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n564), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT85), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n334), .A2(new_n331), .ZN(new_n573));
  OR3_X1    g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n571), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n528), .A2(KEYINPUT26), .A3(new_n492), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n490), .A2(new_n491), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n494), .B2(new_n496), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n523), .A2(new_n527), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n577), .B(KEYINPUT84), .C1(KEYINPUT26), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n523), .ZN(new_n583));
  AND4_X1   g0383(.A1(KEYINPUT26), .A2(new_n492), .A3(new_n523), .A4(new_n527), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n464), .B1(new_n439), .B2(new_n447), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n558), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(new_n500), .A3(new_n532), .A4(new_n528), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n426), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n576), .A2(new_n591), .ZN(G369));
  NOR2_X1   g0392(.A1(new_n467), .A2(new_n533), .ZN(new_n593));
  OR3_X1    g0393(.A1(new_n297), .A2(KEYINPUT27), .A3(G20), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT27), .B1(new_n297), .B2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(G213), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G343), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n593), .B1(new_n448), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n467), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(new_n602));
  INV_X1    g0402(.A(new_n558), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n544), .A2(new_n599), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n561), .B2(new_n604), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G330), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n558), .A2(new_n598), .ZN(new_n611));
  INV_X1    g0411(.A(new_n587), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n593), .A2(new_n611), .B1(new_n612), .B2(new_n599), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n613), .ZN(G399));
  INV_X1    g0414(.A(new_n210), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(G41), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n206), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n517), .A2(G116), .ZN(new_n618));
  INV_X1    g0418(.A(new_n213), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n616), .ZN(new_n620));
  XOR2_X1   g0420(.A(new_n620), .B(KEYINPUT28), .Z(new_n621));
  NAND4_X1  g0421(.A1(new_n489), .A2(new_n510), .A3(new_n462), .A4(new_n555), .ZN(new_n622));
  XOR2_X1   g0422(.A(new_n622), .B(KEYINPUT30), .Z(new_n623));
  NAND3_X1  g0423(.A1(new_n512), .A2(new_n276), .A3(new_n551), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n463), .A2(new_n488), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n598), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT31), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT31), .B(new_n598), .C1(new_n623), .C2(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n562), .A2(new_n599), .B1(new_n632), .B2(KEYINPUT87), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G330), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n467), .A2(new_n603), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n500), .A2(new_n532), .A3(new_n528), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n528), .A2(new_n640), .A3(new_n492), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n641), .B(new_n523), .C1(new_n640), .C2(new_n581), .ZN(new_n642));
  OAI211_X1 g0442(.A(KEYINPUT29), .B(new_n599), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n590), .A2(new_n599), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(KEYINPUT29), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n621), .B1(new_n647), .B2(G1), .ZN(G364));
  NAND2_X1  g0448(.A1(new_n207), .A2(G13), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT88), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G45), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n617), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n608), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(G330), .B2(new_n606), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n207), .A2(G190), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n350), .A2(G179), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(G179), .A2(G200), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(G283), .A2(new_n659), .B1(new_n662), .B2(G329), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT96), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n207), .A2(new_n276), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G200), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n304), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n207), .B1(new_n660), .B2(G190), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(G326), .B1(G294), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT95), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT94), .ZN(new_n672));
  INV_X1    g0472(.A(new_n666), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n304), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n666), .A2(KEYINPUT94), .A3(G190), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(KEYINPUT33), .B(G317), .Z(new_n677));
  OAI211_X1 g0477(.A(new_n664), .B(new_n671), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n276), .A2(G200), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n656), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n258), .B1(new_n681), .B2(G311), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n207), .A2(new_n304), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n657), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n679), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(G303), .A2(new_n685), .B1(new_n687), .B2(G322), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n682), .B(new_n688), .C1(new_n670), .C2(KEYINPUT95), .ZN(new_n689));
  XOR2_X1   g0489(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(KEYINPUT91), .B(G159), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n662), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(G50), .B2(new_n667), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n686), .A2(new_n358), .B1(new_n680), .B2(new_n219), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n658), .A2(new_n221), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n669), .A2(G97), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n693), .A2(new_n691), .A3(new_n662), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n698), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n258), .B1(new_n684), .B2(new_n431), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n244), .B2(new_n676), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n678), .A2(new_n689), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(G20), .B1(KEYINPUT89), .B2(G169), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(KEYINPUT89), .A2(G169), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n215), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT90), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n615), .A2(new_n265), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n712), .A2(G355), .B1(new_n541), .B2(new_n615), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n369), .A2(new_n375), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n210), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n214), .A2(new_n449), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n248), .B2(new_n449), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n713), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n709), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n652), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n710), .B1(new_n711), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n711), .B2(new_n724), .ZN(new_n726));
  INV_X1    g0526(.A(new_n722), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n606), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n655), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(G396));
  INV_X1    g0530(.A(new_n709), .ZN(new_n731));
  INV_X1    g0531(.A(G137), .ZN(new_n732));
  INV_X1    g0532(.A(new_n667), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n676), .A2(new_n310), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT99), .Z(new_n735));
  AOI22_X1  g0535(.A1(new_n681), .A2(new_n693), .B1(new_n687), .B2(G143), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT100), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n658), .A2(new_n244), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(G50), .B2(new_n685), .ZN(new_n742));
  INV_X1    g0542(.A(G132), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n743), .B2(new_n661), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n715), .B(new_n744), .C1(G58), .C2(new_n669), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n699), .B1(new_n733), .B2(new_n548), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n659), .A2(G87), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n541), .B2(new_n680), .ZN(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n686), .A2(new_n750), .B1(new_n661), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n747), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n265), .B1(new_n684), .B2(new_n221), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n753), .B(new_n755), .C1(new_n756), .C2(new_n676), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n731), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n344), .A2(new_n598), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n351), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n353), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n353), .A2(new_n598), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n731), .A2(new_n721), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n766), .A2(new_n721), .B1(G77), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n653), .B1(new_n759), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n644), .B(new_n766), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n636), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n652), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n636), .A2(new_n770), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT101), .Z(G384));
  NOR2_X1   g0575(.A1(new_n650), .A2(new_n206), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n302), .B(new_n598), .C1(new_n279), .C2(new_n565), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n302), .A2(new_n598), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n277), .B1(new_n272), .B2(new_n274), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n307), .B(new_n778), .C1(new_n779), .C2(new_n301), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n766), .ZN(new_n782));
  INV_X1    g0582(.A(new_n632), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n529), .A2(new_n561), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n593), .A2(new_n784), .A3(new_n599), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n596), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n416), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n421), .C1(new_n401), .C2(new_n414), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(KEYINPUT37), .ZN(new_n790));
  INV_X1    g0590(.A(new_n421), .ZN(new_n791));
  INV_X1    g0591(.A(new_n357), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT71), .B1(new_n383), .B2(G68), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n386), .A2(new_n385), .A3(new_n244), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n363), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n285), .B1(new_n795), .B2(new_n399), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n389), .B1(new_n796), .B2(KEYINPUT103), .ZN(new_n797));
  OAI211_X1 g0597(.A(KEYINPUT103), .B(new_n286), .C1(new_n388), .C2(KEYINPUT16), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n792), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n791), .B1(new_n800), .B2(new_n413), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT104), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n399), .B(new_n364), .C1(new_n384), .C2(new_n387), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n286), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT103), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n357), .B1(new_n806), .B2(new_n798), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n802), .B1(new_n807), .B2(new_n596), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n800), .A2(KEYINPUT104), .A3(new_n787), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n801), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n790), .B1(new_n810), .B2(KEYINPUT37), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n425), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT38), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n425), .A2(new_n788), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n789), .B(KEYINPUT37), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT38), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n786), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n810), .A2(KEYINPUT37), .ZN(new_n819));
  INV_X1    g0619(.A(new_n790), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n425), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n809), .A2(new_n808), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(KEYINPUT38), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n783), .A2(new_n785), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT40), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n765), .B1(new_n777), .B2(new_n780), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n818), .A2(KEYINPUT40), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n426), .A2(new_n828), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  INV_X1    g0636(.A(G330), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n821), .B2(new_n824), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT39), .B1(new_n840), .B2(new_n814), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n815), .A2(new_n816), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n813), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT39), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n825), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(KEYINPUT105), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n303), .A2(new_n598), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT105), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n827), .A2(new_n848), .A3(KEYINPUT39), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n781), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n590), .A2(new_n599), .A3(new_n766), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n764), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n855), .A3(new_n764), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n851), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(new_n827), .B1(new_n569), .B2(new_n596), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n426), .B(new_n643), .C1(KEYINPUT29), .C2(new_n645), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n576), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n859), .B(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n776), .B1(new_n839), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n839), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(G116), .A3(new_n216), .A4(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OAI21_X1  g0668(.A(G77), .B1(new_n358), .B2(new_n244), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n243), .B1(new_n869), .B2(new_n213), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(G1), .A3(new_n280), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n864), .A2(new_n868), .A3(new_n871), .ZN(G367));
  OAI21_X1  g0672(.A(new_n500), .B1(new_n497), .B2(new_n599), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n579), .B2(new_n599), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n609), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT107), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n526), .A2(new_n599), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n583), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n580), .B2(new_n877), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT43), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n876), .B(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n492), .B1(new_n874), .B2(new_n467), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n598), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n593), .A2(new_n874), .A3(new_n611), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT106), .Z(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(KEYINPUT42), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(KEYINPUT42), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n879), .A2(KEYINPUT43), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n881), .B(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n616), .B(KEYINPUT41), .Z(new_n891));
  NAND2_X1  g0691(.A1(new_n593), .A2(new_n611), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n602), .B2(new_n611), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(new_n608), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n647), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n613), .A2(new_n874), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT45), .Z(new_n898));
  NOR2_X1   g0698(.A1(new_n613), .A2(new_n874), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT44), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(new_n610), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n891), .B1(new_n904), .B2(new_n647), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n651), .A2(G1), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n723), .B1(new_n210), .B2(new_n341), .C1(new_n238), .C2(new_n716), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n653), .ZN(new_n909));
  INV_X1    g0709(.A(new_n676), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n714), .B1(new_n910), .B2(G294), .ZN(new_n911));
  AOI22_X1  g0711(.A1(G303), .A2(new_n687), .B1(new_n662), .B2(G317), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n468), .B2(new_n658), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n685), .A2(KEYINPUT46), .A3(G116), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n733), .B2(new_n751), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT46), .B1(new_n685), .B2(G116), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n680), .A2(new_n756), .B1(new_n668), .B2(new_n221), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT109), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n910), .A2(new_n693), .B1(G50), .B2(new_n681), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT110), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n661), .A2(new_n732), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n658), .A2(new_n219), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(G150), .C2(new_n687), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n668), .A2(new_n244), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n258), .B1(new_n684), .B2(new_n358), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n927), .B(new_n928), .C1(G143), .C2(new_n667), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n923), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n920), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT47), .Z(new_n933));
  OAI221_X1 g0733(.A(new_n909), .B1(new_n879), .B2(new_n727), .C1(new_n731), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n907), .A2(new_n934), .ZN(G387));
  OR2_X1    g0735(.A1(new_n602), .A2(new_n727), .ZN(new_n936));
  INV_X1    g0736(.A(new_n712), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n937), .A2(new_n618), .B1(G107), .B2(new_n210), .ZN(new_n938));
  INV_X1    g0738(.A(new_n234), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n716), .B1(new_n939), .B2(G45), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n618), .B(new_n449), .C1(new_n244), .C2(new_n219), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT50), .B1(new_n309), .B2(G50), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n309), .A2(KEYINPUT50), .A3(G50), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n938), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n723), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n653), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n684), .A2(new_n750), .B1(new_n668), .B2(new_n756), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G317), .A2(new_n687), .B1(new_n681), .B2(G303), .ZN(new_n951));
  INV_X1    g0751(.A(G322), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n952), .B2(new_n733), .C1(new_n676), .C2(new_n751), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT48), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT49), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G116), .A2(new_n659), .B1(new_n662), .B2(G326), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n715), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT114), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n956), .B2(new_n957), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n685), .A2(G77), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n310), .B2(new_n661), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n964), .A2(KEYINPUT112), .B1(G97), .B2(new_n659), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n965), .B(new_n714), .C1(KEYINPUT112), .C2(new_n964), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT113), .Z(new_n967));
  OAI22_X1  g0767(.A1(new_n686), .A2(new_n202), .B1(new_n680), .B2(new_n244), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n341), .A2(new_n668), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G159), .C2(new_n667), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n309), .B2(new_n676), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n958), .A2(new_n962), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n949), .B1(new_n972), .B2(new_n709), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n894), .A2(new_n906), .B1(new_n936), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n895), .A2(new_n616), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n894), .A2(new_n647), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G393));
  AND2_X1   g0777(.A1(new_n894), .A2(new_n647), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n904), .B(new_n616), .C1(new_n978), .C2(new_n902), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n902), .A2(new_n906), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n723), .B1(new_n468), .B2(new_n210), .C1(new_n716), .C2(new_n242), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n653), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n668), .A2(new_n219), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n337), .B2(new_n681), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n676), .B2(new_n202), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT115), .Z(new_n986));
  AOI22_X1  g0786(.A1(new_n667), .A2(G150), .B1(new_n687), .B2(G159), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT51), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n748), .B1(new_n244), .B2(new_n684), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n989), .B(new_n715), .C1(G143), .C2(new_n662), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT116), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n667), .A2(G317), .B1(new_n687), .B2(G311), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT52), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n910), .A2(G303), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n680), .A2(new_n750), .B1(new_n661), .B2(new_n952), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G283), .B2(new_n685), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n258), .B(new_n697), .C1(G116), .C2(new_n669), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n991), .A2(new_n992), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n993), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n982), .B1(new_n1002), .B2(new_n709), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n874), .B2(new_n727), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n979), .A2(new_n980), .A3(new_n1004), .ZN(G390));
  NOR2_X1   g0805(.A1(new_n765), .A2(new_n837), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n828), .A2(new_n781), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n854), .A2(new_n856), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n847), .B1(new_n1009), .B2(new_n781), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n846), .B2(new_n849), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n599), .B(new_n762), .C1(new_n639), .C2(new_n642), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n764), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n847), .B1(new_n1013), .B2(new_n781), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n825), .A2(new_n843), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1008), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1006), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n633), .B2(new_n634), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n781), .ZN(new_n1021));
  AOI211_X1 g0821(.A(KEYINPUT105), .B(new_n844), .C1(new_n825), .C2(new_n826), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n848), .B1(new_n827), .B2(KEYINPUT39), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n845), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1016), .B(new_n1021), .C1(new_n1024), .C2(new_n1010), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1007), .B1(new_n1020), .B2(new_n781), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n781), .B1(new_n828), .B2(new_n1006), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n1013), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1027), .A2(new_n1009), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n828), .A2(G330), .A3(new_n425), .A4(new_n355), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT117), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n426), .A2(KEYINPUT117), .A3(G330), .A4(new_n828), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n576), .A3(new_n860), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1026), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1018), .A2(new_n1025), .A3(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n616), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1018), .A2(new_n1025), .A3(new_n906), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n653), .B1(new_n337), .B2(new_n767), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT118), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n680), .A2(new_n468), .B1(new_n661), .B2(new_n750), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n741), .B(new_n1045), .C1(G116), .C2(new_n687), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n265), .B1(new_n684), .B2(new_n431), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n983), .B(new_n1047), .C1(G283), .C2(new_n667), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n221), .C2(new_n676), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n685), .A2(G150), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT53), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G159), .B2(new_n669), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT54), .B(G143), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n687), .A2(G132), .B1(new_n681), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(G128), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n733), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1052), .B(new_n1058), .C1(new_n732), .C2(new_n676), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n258), .B1(new_n658), .B2(new_n202), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G125), .B2(new_n662), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT119), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1049), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1044), .B1(new_n1063), .B2(new_n709), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1024), .B2(new_n721), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1041), .A2(new_n1042), .A3(new_n1065), .ZN(G378));
  INV_X1    g0866(.A(new_n1036), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1040), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n332), .A2(new_n787), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n335), .B(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n832), .B2(new_n837), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n829), .B1(new_n1015), .B2(new_n786), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n825), .B2(new_n826), .ZN(new_n1077));
  OAI211_X1 g0877(.A(G330), .B(new_n1072), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n859), .A3(KEYINPUT123), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n859), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT123), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1074), .A2(new_n850), .A3(new_n1078), .A4(new_n858), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1068), .A2(KEYINPUT57), .A3(new_n1080), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT124), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1079), .A2(new_n859), .A3(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT122), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1081), .A2(new_n1088), .A3(new_n1083), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1068), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT57), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1040), .B2(new_n1067), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT124), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1080), .A4(new_n1084), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1086), .A2(new_n1092), .A3(new_n616), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1089), .A2(new_n906), .A3(new_n1087), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n653), .B1(G50), .B2(new_n767), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n715), .B1(new_n676), .B2(new_n468), .ZN(new_n1099));
  AOI21_X1  g0899(.A(G41), .B1(new_n685), .B2(G77), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n244), .B2(new_n668), .C1(new_n733), .C2(new_n541), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n341), .A2(new_n680), .B1(new_n358), .B2(new_n658), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n686), .A2(new_n221), .B1(new_n661), .B2(new_n756), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT58), .Z(new_n1105));
  AOI21_X1  g0905(.A(G41), .B1(new_n714), .B2(G33), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1056), .A2(new_n686), .B1(new_n684), .B2(new_n1053), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G137), .B2(new_n681), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n667), .A2(G125), .B1(G150), .B2(new_n669), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n676), .C2(new_n743), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT59), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n662), .A2(G124), .ZN(new_n1113));
  AOI211_X1 g0913(.A(G33), .B(G41), .C1(new_n693), .C2(new_n659), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1105), .B1(G50), .B2(new_n1106), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT121), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n731), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1098), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n1072), .B2(new_n721), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1096), .A2(new_n1123), .ZN(G375));
  NOR2_X1   g0924(.A1(new_n1037), .A2(new_n891), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1030), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n851), .A2(new_n720), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n653), .B1(G68), .B2(new_n767), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n681), .B1(new_n662), .B2(G303), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n468), .B2(new_n684), .C1(new_n756), .C2(new_n686), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n969), .B(new_n1132), .C1(G294), .C2(new_n667), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n925), .A2(new_n258), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT125), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(new_n541), .C2(new_n676), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n715), .B1(new_n910), .B2(new_n1054), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n680), .A2(new_n310), .B1(new_n661), .B2(new_n1056), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G137), .B2(new_n687), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n668), .A2(new_n202), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n684), .A2(new_n361), .B1(new_n658), .B2(new_n358), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(G132), .C2(new_n667), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1136), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1130), .B1(new_n1144), .B2(new_n709), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1128), .A2(new_n906), .B1(new_n1129), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1127), .A2(new_n1146), .ZN(G381));
  INV_X1    g0947(.A(G390), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1148), .A2(new_n1146), .A3(new_n1127), .A4(new_n1149), .ZN(new_n1150));
  OR4_X1    g0950(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1150), .ZN(G407));
  INV_X1    g0951(.A(G378), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n597), .A2(G213), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G407), .B(G213), .C1(G375), .C2(new_n1155), .ZN(G409));
  INV_X1    g0956(.A(KEYINPUT61), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1096), .A2(G378), .A3(new_n1123), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1090), .A2(new_n891), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1084), .A2(new_n906), .A3(new_n1080), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1122), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1152), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n616), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT60), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n1126), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT126), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1030), .A2(new_n1036), .A3(KEYINPUT60), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1146), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G384), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G384), .B(new_n1146), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1153), .A2(KEYINPUT127), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1154), .A2(G2897), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .A4(new_n1175), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1157), .B1(new_n1163), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT63), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1153), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(G393), .B(new_n729), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(G387), .A2(new_n1148), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G387), .A2(new_n1148), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1190), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1187), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1163), .A2(KEYINPUT63), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1183), .A2(new_n1188), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT62), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1163), .A2(new_n1202), .A3(new_n1199), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1163), .B2(new_n1199), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1203), .A2(new_n1182), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1201), .B1(new_n1205), .B2(new_n1198), .ZN(G405));
  NAND2_X1  g1006(.A1(G375), .A2(new_n1152), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1158), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1199), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1187), .A3(new_n1158), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(new_n1197), .ZN(G402));
endmodule


