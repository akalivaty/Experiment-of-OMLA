//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(KEYINPUT66), .ZN(new_n243));
  AND2_X1   g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n243), .B1(new_n244), .B2(new_n209), .ZN(new_n245));
  AND2_X1   g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(KEYINPUT66), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n244), .A2(new_n209), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G223), .A3(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n255), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n253), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n245), .A2(new_n252), .A3(new_n248), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n245), .A2(new_n248), .A3(new_n264), .A4(new_n252), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n209), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G150), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n210), .A2(G33), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n210), .B1(new_n201), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n272), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n278), .B1(new_n251), .B2(G20), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(new_n284), .B1(new_n278), .B2(new_n282), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n261), .A2(new_n267), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n270), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(G200), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(KEYINPUT68), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n286), .B(KEYINPUT9), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n261), .A2(new_n267), .A3(G190), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n295), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G33), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n300), .A2(new_n302), .A3(G226), .A4(new_n256), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n300), .A2(new_n302), .A3(G232), .A4(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n254), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n244), .A2(new_n243), .A3(new_n209), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT66), .B1(new_n246), .B2(new_n247), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n252), .A2(new_n250), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n266), .A2(G238), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n216), .B1(new_n263), .B2(new_n265), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT13), .B1(new_n318), .B2(new_n313), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(new_n273), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n322), .A2(new_n278), .B1(new_n210), .B2(G68), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n276), .A2(new_n259), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n272), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n281), .A2(G68), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n328), .C2(new_n327), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n251), .A2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n283), .A2(G68), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n321), .B(new_n336), .C1(new_n337), .C2(new_n320), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G107), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(new_n341), .C2(new_n255), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n254), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n312), .ZN(new_n344));
  INV_X1    g0144(.A(G244), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n263), .B2(new_n265), .ZN(new_n346));
  OAI21_X1  g0146(.A(G200), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n253), .B1(new_n254), .B2(new_n342), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n266), .A2(G244), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G190), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n275), .A2(new_n322), .B1(new_n210), .B2(new_n259), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n276), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n272), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n333), .A2(G77), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n283), .A2(new_n356), .B1(new_n259), .B2(new_n282), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n347), .A2(new_n350), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n269), .B1(new_n344), .B2(new_n346), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n357), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n348), .A2(new_n349), .A3(new_n287), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n338), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n298), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n318), .A2(new_n313), .A3(KEYINPUT13), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n320), .B2(G169), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n335), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  AND2_X1   g0174(.A1(G226), .A2(G1698), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n255), .B2(new_n375), .ZN(new_n376));
  AND4_X1   g0176(.A1(new_n374), .A2(new_n300), .A3(new_n302), .A4(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n255), .A2(G223), .A3(new_n256), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT74), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n300), .A2(new_n302), .A3(new_n375), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT73), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n255), .A2(new_n374), .A3(new_n375), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n380), .A4(new_n379), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n254), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n312), .B1(new_n390), .B2(new_n262), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(G179), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n254), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n380), .B(new_n379), .C1(new_n376), .C2(new_n377), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(KEYINPUT74), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n391), .B1(new_n396), .B2(new_n388), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(new_n269), .ZN(new_n398));
  INV_X1    g0198(.A(new_n283), .ZN(new_n399));
  INV_X1    g0199(.A(new_n275), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n333), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n399), .A2(new_n401), .B1(new_n281), .B2(new_n400), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n273), .A2(G159), .ZN(new_n405));
  AND2_X1   g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(KEYINPUT70), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT70), .ZN(new_n409));
  XNOR2_X1  g0209(.A(G58), .B(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n404), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n409), .A3(G20), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT71), .A4(new_n405), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n300), .A2(new_n302), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n418), .B2(new_n210), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n255), .B2(G20), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT72), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G68), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT16), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n423), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(G68), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n412), .A2(new_n415), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n272), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n403), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n398), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  AOI211_X1 g0236(.A(G190), .B(new_n391), .C1(new_n396), .C2(new_n388), .ZN(new_n437));
  AOI21_X1  g0237(.A(G200), .B1(new_n389), .B2(new_n392), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n439), .B2(new_n433), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n398), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n389), .A2(new_n337), .A3(new_n392), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n397), .B2(G200), .ZN(new_n444));
  INV_X1    g0244(.A(new_n272), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n416), .B2(new_n429), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n420), .B(G20), .C1(new_n300), .C2(new_n302), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n417), .B1(new_n419), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT72), .B1(new_n422), .B2(KEYINPUT7), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n215), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n427), .B1(new_n450), .B2(new_n431), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n402), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n444), .A2(new_n452), .A3(KEYINPUT17), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n435), .A2(new_n440), .A3(new_n442), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n365), .A2(new_n373), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT75), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n365), .A2(new_n455), .A3(new_n458), .A4(new_n373), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n251), .A2(G33), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n283), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n282), .A2(KEYINPUT25), .A3(new_n341), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT25), .B1(new_n282), .B2(new_n341), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n462), .A2(new_n341), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n255), .A2(new_n466), .A3(new_n210), .A4(G87), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n300), .A2(new_n302), .A3(new_n210), .A4(G87), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT81), .B(KEYINPUT22), .Z(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n210), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n341), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n299), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n472), .A2(new_n473), .B1(new_n475), .B2(new_n210), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n467), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n478), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n467), .A2(new_n470), .A3(new_n476), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n465), .B1(new_n482), .B2(new_n272), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n488), .A2(new_n245), .A3(new_n248), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n300), .A2(new_n302), .A3(G257), .A4(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n300), .A2(new_n302), .A3(G250), .A4(new_n256), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT83), .B(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n299), .C2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(G264), .A2(new_n489), .B1(new_n493), .B2(new_n254), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n485), .B(G274), .C1(new_n487), .C2(new_n486), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n310), .A2(new_n496), .A3(KEYINPUT77), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT77), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n249), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n494), .A2(new_n287), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(G169), .B1(new_n494), .B2(new_n500), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n483), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n494), .A2(KEYINPUT84), .A3(new_n500), .A4(new_n337), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(new_n500), .ZN(new_n506));
  INV_X1    g0306(.A(G200), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n506), .A2(G190), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n510), .B2(new_n483), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n300), .A2(new_n302), .A3(G244), .A4(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n300), .A2(new_n302), .A3(G238), .A4(new_n256), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n299), .C2(new_n474), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n254), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n485), .A2(G250), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n484), .A2(G1), .A3(G274), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n310), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n352), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n281), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n255), .A2(new_n210), .A3(G68), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n276), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n217), .A2(new_n526), .A3(new_n341), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT78), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n217), .A3(new_n526), .A4(new_n341), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n533), .A2(new_n210), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n524), .B(new_n527), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n523), .B1(new_n535), .B2(new_n272), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n283), .A2(new_n461), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(KEYINPUT79), .A3(G87), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n462), .B2(new_n217), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n514), .A2(new_n254), .B1(new_n310), .B2(new_n518), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n521), .A2(new_n536), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(new_n522), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n524), .A2(new_n527), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n534), .B1(new_n529), .B2(new_n531), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n272), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n523), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n287), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(G169), .C2(new_n542), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n341), .B1(new_n448), .B2(new_n449), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n526), .A2(new_n341), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n341), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G20), .B1(G77), .B2(new_n273), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n272), .B1(new_n554), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT76), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n462), .A2(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n281), .A2(new_n526), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n564), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n300), .A2(new_n302), .A3(G250), .A4(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G283), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n300), .A2(new_n302), .A3(G244), .A4(new_n256), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n254), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n489), .A2(G257), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n500), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n497), .A2(new_n499), .B1(new_n489), .B2(G257), .ZN(new_n581));
  AOI21_X1  g0381(.A(G200), .B1(new_n581), .B2(new_n577), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n563), .B(new_n570), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n269), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n287), .A3(new_n577), .ZN(new_n585));
  INV_X1    g0385(.A(new_n569), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n567), .ZN(new_n587));
  OAI21_X1  g0387(.A(G107), .B1(new_n421), .B2(new_n424), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n445), .B1(new_n588), .B2(new_n561), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n584), .B(new_n585), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n553), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n281), .A2(G116), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n537), .B2(G116), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n271), .A2(new_n209), .B1(G20), .B2(new_n474), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n572), .B(new_n210), .C1(G33), .C2(new_n526), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(KEYINPUT80), .A3(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g0397(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n594), .B2(new_n595), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n489), .A2(G270), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n300), .A2(new_n302), .A3(G264), .A4(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n300), .A2(new_n302), .A3(G257), .A4(new_n256), .ZN(new_n604));
  INV_X1    g0404(.A(G303), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n255), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n254), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT77), .B1(new_n310), .B2(new_n496), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n249), .A2(new_n495), .A3(new_n498), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n602), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n610), .A3(G169), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n601), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(G200), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n337), .C2(new_n610), .ZN(new_n616));
  INV_X1    g0416(.A(new_n610), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(G179), .A3(new_n601), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n601), .A2(new_n610), .A3(KEYINPUT21), .A4(G169), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n613), .A2(new_n616), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n460), .A2(new_n511), .A3(new_n591), .A4(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n442), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n441), .B1(new_n398), .B2(new_n433), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n362), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n338), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n373), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(KEYINPUT85), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n440), .A2(new_n453), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n627), .B2(KEYINPUT85), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n292), .B(new_n295), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n289), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n483), .A2(new_n501), .A3(new_n502), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n618), .A2(new_n619), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n613), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n510), .A2(new_n483), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n591), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n590), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .A3(new_n553), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n544), .A2(new_n552), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n590), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n552), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n460), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n635), .A2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n637), .A2(new_n613), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n251), .A2(new_n210), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n614), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n620), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n659), .B(KEYINPUT86), .C1(new_n660), .C2(new_n658), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G330), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n511), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n483), .A2(new_n657), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT87), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n503), .B2(new_n656), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n650), .A2(new_n657), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n671), .A2(new_n676), .B1(new_n503), .B2(new_n657), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(G399));
  NAND2_X1  g0478(.A1(new_n532), .A2(new_n474), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n206), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n213), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n647), .A2(new_n657), .ZN(new_n687));
  XNOR2_X1  g0487(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n642), .A2(KEYINPUT91), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n642), .A2(KEYINPUT91), .A3(new_n645), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n640), .A3(new_n552), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n617), .A2(G179), .A3(new_n577), .A4(new_n581), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n493), .A2(new_n254), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n310), .A2(G264), .A3(new_n488), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n515), .A3(new_n698), .A4(new_n519), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT88), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT88), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n494), .A2(new_n542), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n695), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n579), .A2(new_n610), .A3(new_n287), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n702), .A4(new_n700), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n542), .B(KEYINPUT89), .ZN(new_n707));
  AOI21_X1  g0507(.A(G179), .B1(new_n581), .B2(new_n577), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n506), .A3(new_n610), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n656), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n591), .A2(new_n511), .A3(new_n620), .A4(new_n657), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n694), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n686), .B1(new_n718), .B2(G1), .ZN(G364));
  NAND2_X1  g0519(.A1(new_n663), .A2(new_n664), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  AND2_X1   g0521(.A1(new_n210), .A2(G13), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n251), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n721), .B(new_n666), .C1(new_n682), .C2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n663), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n210), .A2(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G190), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G87), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G159), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n738));
  OAI21_X1  g0538(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n210), .A2(new_n287), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n337), .A3(G200), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n255), .B1(new_n741), .B2(new_n215), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n734), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(G77), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n730), .A2(new_n337), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n341), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n740), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n507), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G50), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n210), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n748), .A2(G200), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G97), .A2(new_n753), .B1(new_n754), .B2(G58), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n745), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n739), .B(new_n756), .C1(new_n737), .C2(new_n738), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n759));
  INV_X1    g0559(.A(new_n754), .ZN(new_n760));
  INV_X1    g0560(.A(G322), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(new_n605), .B2(new_n731), .ZN(new_n762));
  INV_X1    g0562(.A(new_n746), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G283), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  INV_X1    g0565(.A(G329), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n741), .A2(new_n765), .B1(new_n766), .B2(new_n735), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n255), .B(new_n767), .C1(G311), .C2(new_n744), .ZN(new_n768));
  INV_X1    g0568(.A(new_n492), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(new_n753), .B1(new_n749), .B2(G326), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n758), .A2(new_n759), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n209), .B1(G20), .B2(new_n269), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n682), .B(new_n724), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n238), .A2(new_n484), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n681), .A2(new_n255), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n213), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n776), .B2(new_n775), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n681), .A2(new_n418), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G355), .B1(new_n474), .B2(new_n681), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT95), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(KEYINPUT95), .A3(new_n784), .ZN(new_n786));
  INV_X1    g0586(.A(new_n728), .ZN(new_n787));
  INV_X1    g0587(.A(new_n773), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n729), .B(new_n774), .C1(new_n785), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n725), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  INV_X1    g0594(.A(new_n741), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G150), .B1(new_n744), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(new_n749), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  INV_X1    g0598(.A(G143), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(new_n797), .B2(new_n798), .C1(new_n799), .C2(new_n760), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  INV_X1    g0604(.A(G58), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n255), .B1(new_n735), .B2(new_n804), .C1(new_n752), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n763), .A2(G68), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n278), .B2(new_n731), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n802), .A2(new_n803), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n760), .A2(new_n810), .B1(new_n217), .B2(new_n746), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n741), .A2(new_n812), .B1(new_n743), .B2(new_n474), .ZN(new_n813));
  INV_X1    g0613(.A(new_n735), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n255), .B(new_n813), .C1(G311), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G97), .A2(new_n753), .B1(new_n749), .B2(G303), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n811), .B(new_n817), .C1(G107), .C2(new_n732), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n773), .B1(new_n809), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n724), .A2(new_n682), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n773), .A2(new_n726), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT99), .Z(new_n822));
  OAI211_X1 g0622(.A(new_n819), .B(new_n820), .C1(G77), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n360), .A2(new_n656), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n358), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n362), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n625), .A2(new_n657), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n823), .B1(new_n832), .B2(new_n726), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n687), .B1(new_n830), .B2(new_n829), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n647), .A3(new_n657), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n717), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n820), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n717), .A3(new_n835), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  AOI211_X1 g0640(.A(new_n474), .B(new_n212), .C1(new_n560), .C2(KEYINPUT35), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(KEYINPUT35), .B2(new_n560), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT36), .Z(new_n843));
  OR3_X1    g0643(.A1(new_n213), .A2(new_n259), .A3(new_n406), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n278), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n251), .B(G13), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT103), .B1(new_n694), .B2(new_n460), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n694), .A2(KEYINPUT103), .A3(new_n460), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n634), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT104), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n428), .A2(G68), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n416), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n403), .B1(new_n855), .B2(new_n432), .ZN(new_n856));
  INV_X1    g0656(.A(new_n654), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n454), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n398), .A2(new_n856), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n444), .A2(new_n452), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n287), .B(new_n391), .C1(new_n396), .C2(new_n388), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n269), .B1(new_n389), .B2(new_n392), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT102), .B1(new_n867), .B2(new_n452), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n433), .A2(new_n857), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT37), .B1(new_n444), .B2(new_n452), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n398), .A2(new_n433), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n860), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n454), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n434), .A2(new_n862), .A3(new_n869), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n873), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n853), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n858), .B1(new_n629), .B2(new_n624), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n398), .A2(new_n433), .A3(new_n871), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n871), .B1(new_n398), .B2(new_n433), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n862), .A2(new_n869), .A3(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n887), .A2(new_n889), .B1(KEYINPUT37), .B2(new_n863), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n883), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n860), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n373), .A2(KEYINPUT101), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n335), .C1(new_n371), .C2(new_n372), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n656), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n882), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n335), .A2(new_n656), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n338), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n371), .A2(new_n372), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n338), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n335), .A3(new_n656), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n828), .B2(new_n835), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n891), .A2(new_n892), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n654), .B1(new_n622), .B2(new_n623), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n899), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n852), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n716), .A2(new_n831), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n869), .B1(new_n629), .B2(new_n624), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n887), .A2(new_n889), .B1(KEYINPUT37), .B2(new_n878), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n883), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n919), .B2(new_n892), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n915), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n460), .A2(new_n716), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n664), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n912), .A2(KEYINPUT105), .A3(new_n924), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n251), .B2(new_n722), .C1(new_n912), .C2(new_n924), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT105), .B1(new_n912), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n847), .B1(new_n926), .B2(new_n927), .ZN(G367));
  NOR3_X1   g0728(.A1(new_n234), .A2(new_n681), .A3(new_n255), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n790), .B1(new_n206), .B2(new_n352), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n820), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n797), .A2(new_n799), .B1(new_n731), .B2(new_n805), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(G68), .B2(new_n753), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n418), .B1(new_n814), .B2(G137), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n795), .A2(G159), .B1(new_n744), .B2(G50), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n754), .A2(G150), .B1(new_n763), .B2(G77), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n731), .A2(new_n474), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT46), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G107), .A2(new_n753), .B1(new_n749), .B2(G311), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n754), .A2(G303), .B1(new_n763), .B2(G97), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n255), .B1(new_n744), .B2(G283), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT110), .B(G317), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n795), .A2(new_n769), .B1(new_n814), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n940), .A2(new_n941), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n937), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n931), .B1(new_n947), .B2(new_n773), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n536), .A2(new_n541), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n656), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n553), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n552), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n948), .B1(new_n787), .B2(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n675), .B1(new_n636), .B2(new_n657), .C1(new_n667), .C2(new_n670), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n671), .A2(new_n676), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n665), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n666), .A2(new_n957), .A3(new_n956), .A4(new_n958), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n718), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(new_n677), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n641), .A2(new_n656), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n656), .B1(new_n587), .B2(new_n589), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n583), .A2(new_n590), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT106), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n967), .A2(KEYINPUT106), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n965), .B1(new_n966), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n677), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n677), .B2(new_n974), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n966), .A2(new_n975), .A3(KEYINPUT44), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(KEYINPUT108), .A3(new_n980), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n674), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n978), .A2(new_n981), .ZN(new_n986));
  INV_X1    g0786(.A(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n673), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n964), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n718), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n682), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n724), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n975), .A2(new_n957), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT42), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n641), .B1(new_n974), .B2(new_n503), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n656), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n997), .B2(new_n996), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n995), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n953), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT43), .B2(new_n953), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n953), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n995), .A2(new_n999), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n674), .A2(new_n975), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1001), .A2(new_n1006), .A3(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n954), .B1(new_n993), .B2(new_n1010), .ZN(G387));
  AOI21_X1  g0811(.A(new_n255), .B1(new_n814), .B2(G326), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n474), .B2(new_n746), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n795), .A2(G311), .B1(new_n744), .B2(G303), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n761), .B2(new_n797), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n754), .B2(new_n943), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT112), .Z(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n753), .A2(G283), .B1(new_n732), .B2(new_n769), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT49), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G68), .A2(new_n744), .B1(new_n814), .B2(G150), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1026), .B(new_n255), .C1(new_n275), .C2(new_n741), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n753), .A2(new_n522), .B1(new_n732), .B2(G77), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n278), .B2(new_n760), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n797), .A2(new_n736), .B1(new_n746), .B2(new_n526), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n773), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n275), .A2(G50), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g0834(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1035), .C1(new_n1036), .C2(new_n679), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n680), .A2(KEYINPUT111), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n778), .B1(new_n1037), .B2(new_n1038), .C1(new_n484), .C2(new_n230), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n679), .A2(new_n783), .B1(new_n341), .B2(new_n681), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n790), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1032), .A2(new_n820), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n672), .B2(new_n728), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n724), .B2(new_n962), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n962), .A2(new_n718), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n963), .A2(new_n682), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n985), .A2(new_n988), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n963), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n682), .A3(new_n989), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n985), .A2(new_n724), .A3(new_n988), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n790), .B1(new_n526), .B2(new_n206), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n241), .A2(new_n778), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n820), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n418), .B1(new_n814), .B2(G143), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n215), .B2(new_n731), .C1(new_n217), .C2(new_n746), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT114), .Z(new_n1059));
  AOI22_X1  g0859(.A1(G150), .A2(new_n749), .B1(new_n754), .B2(G159), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n752), .A2(new_n259), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n741), .A2(new_n278), .B1(new_n743), .B2(new_n275), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n418), .B1(new_n735), .B2(new_n761), .C1(new_n810), .C2(new_n743), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n747), .B(new_n1065), .C1(G283), .C2(new_n732), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n753), .A2(G116), .B1(new_n795), .B2(G303), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT115), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G311), .A2(new_n754), .B1(new_n749), .B2(G317), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT52), .Z(new_n1073));
  AOI22_X1  g0873(.A1(new_n1059), .A2(new_n1064), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1056), .B1(new_n788), .B2(new_n1074), .C1(new_n974), .C2(new_n787), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1051), .A2(new_n1052), .A3(new_n1075), .ZN(G390));
  NOR2_X1   g0876(.A1(new_n913), .A2(new_n664), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n902), .A2(new_n905), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n692), .A2(new_n657), .A3(new_n831), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1080), .A2(new_n828), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n906), .B1(new_n913), .B2(new_n664), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1079), .A2(new_n1082), .B1(new_n828), .B2(new_n835), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n460), .A2(new_n717), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n851), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n835), .A2(new_n828), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1078), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n898), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1090), .A2(new_n1091), .B1(new_n882), .B2(new_n893), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n906), .B1(new_n1080), .B2(new_n828), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n875), .A2(new_n881), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n898), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1078), .B(new_n1077), .C1(new_n1092), .C2(new_n1095), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1093), .A2(new_n898), .A3(new_n1094), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n882), .A2(new_n893), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n907), .B2(new_n898), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1099), .A3(new_n1079), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n683), .B1(new_n1088), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1101), .B2(new_n1088), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(new_n726), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n820), .B1(new_n822), .B2(new_n400), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n743), .A2(new_n526), .B1(new_n735), .B2(new_n810), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n255), .B(new_n1107), .C1(G107), .C2(new_n795), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n733), .A3(new_n807), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1062), .B1(G283), .B2(new_n749), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n474), .B2(new_n760), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n732), .A2(G150), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n255), .B1(new_n741), .B2(new_n798), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G125), .B2(new_n814), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G159), .A2(new_n753), .B1(new_n749), .B2(G128), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT116), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n744), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n754), .A2(G132), .B1(new_n763), .B2(G50), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1109), .A2(new_n1111), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1106), .B1(new_n1122), .B2(new_n773), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1104), .A2(new_n724), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1103), .A2(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(new_n821), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n820), .B1(G50), .B2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n760), .A2(new_n341), .B1(new_n805), .B2(new_n746), .ZN(new_n1128));
  INV_X1    g0928(.A(G41), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n418), .A2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n741), .A2(new_n526), .B1(new_n735), .B2(new_n812), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n522), .C2(new_n744), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n215), .B2(new_n752), .C1(new_n259), .C2(new_n731), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1128), .B(new_n1133), .C1(G116), .C2(new_n749), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT58), .Z(new_n1135));
  OAI211_X1 g0935(.A(new_n1130), .B(new_n278), .C1(G33), .C2(G41), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n741), .A2(new_n804), .B1(new_n743), .B2(new_n798), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G150), .B2(new_n753), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G125), .A2(new_n749), .B1(new_n754), .B2(G128), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1118), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1139), .C1(new_n731), .C2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1143));
  OR2_X1    g0943(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n814), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1146), .A2(new_n299), .A3(new_n1129), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1143), .B(new_n1147), .C1(new_n736), .C2(new_n746), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1135), .B(new_n1136), .C1(new_n1142), .C2(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n788), .B1(new_n1149), .B2(KEYINPUT118), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1127), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n298), .A2(new_n286), .A3(new_n857), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n286), .A2(new_n857), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n632), .A2(new_n289), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n726), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1159), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT40), .B1(new_n875), .B2(new_n881), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1078), .A2(new_n716), .A3(new_n831), .ZN(new_n1165));
  OAI21_X1  g0965(.A(G330), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1163), .B1(new_n1166), .B2(new_n915), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n664), .B1(new_n920), .B2(new_n914), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT38), .B1(new_n860), .B2(new_n874), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n875), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n916), .B1(new_n1170), .B2(new_n1165), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1171), .A3(new_n1159), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1172), .A3(new_n911), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT120), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1167), .A2(new_n1172), .A3(new_n1175), .A4(new_n911), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n911), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT119), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1162), .B1(new_n1184), .B2(new_n724), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n851), .B(new_n1087), .C1(new_n1101), .C2(new_n1085), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n694), .A2(KEYINPUT103), .A3(new_n460), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n635), .B(new_n1087), .C1(new_n1188), .C2(new_n848), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1104), .B2(new_n1086), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1173), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n911), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n682), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1187), .B2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1085), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT121), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n992), .A3(new_n1088), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n820), .B1(new_n822), .B2(G68), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n744), .A2(G150), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n418), .B(new_n1200), .C1(G128), .C2(new_n814), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n749), .A2(G132), .B1(new_n763), .B2(G58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n1140), .C2(new_n741), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n753), .A2(G50), .B1(new_n732), .B2(G159), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n798), .B2(new_n760), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n418), .B1(new_n746), .B2(new_n259), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT122), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n743), .A2(new_n341), .B1(new_n735), .B2(new_n605), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G116), .B2(new_n795), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G283), .A2(new_n754), .B1(new_n749), .B2(G294), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n753), .A2(new_n522), .B1(new_n732), .B2(G97), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1203), .A2(new_n1205), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1199), .B1(new_n1213), .B2(new_n773), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1078), .B2(new_n727), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1085), .B2(new_n723), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1198), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G387), .ZN(new_n1219));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  OR4_X1    g1022(.A1(G378), .A2(G375), .A3(new_n1222), .A4(G381), .ZN(G407));
  INV_X1    g1023(.A(G378), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n655), .A2(G213), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G375), .C2(new_n1227), .ZN(G409));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1220), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(G393), .B(new_n793), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G390), .B(new_n954), .C1(new_n993), .C2(new_n1010), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1185), .C1(new_n1187), .C2(new_n1194), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n724), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1180), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT119), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1174), .A2(new_n1176), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1186), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1161), .B(new_n1238), .C1(new_n1243), .C2(new_n991), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1224), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1226), .B1(new_n1237), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n682), .B1(new_n1196), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1088), .A2(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1197), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n839), .B1(new_n1251), .B2(new_n1216), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1196), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT121), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1196), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1249), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(G384), .A3(new_n1217), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1247), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1236), .B1(new_n1262), .B2(KEYINPUT63), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1226), .A2(G2897), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1225), .A2(KEYINPUT124), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1265), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1261), .A2(new_n1270), .A3(new_n1267), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1264), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1263), .B(new_n1274), .C1(KEYINPUT63), .C2(new_n1262), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1247), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT62), .B1(new_n1247), .B2(new_n1261), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1246), .A2(new_n1278), .A3(new_n1266), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1235), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1234), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(KEYINPUT57), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1194), .B1(new_n1243), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n724), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1161), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1224), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1237), .A3(new_n1261), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1288), .A2(new_n1237), .A3(new_n1261), .A4(KEYINPUT125), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1261), .B1(new_n1288), .B2(new_n1237), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1234), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1281), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1234), .A2(new_n1294), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1293), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT126), .B1(new_n1293), .B2(new_n1302), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1301), .A2(new_n1305), .ZN(G402));
endmodule


