//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(G20), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G50), .B(G68), .Z(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G41), .ZN(new_n243));
  INV_X1    g0043(.A(G45), .ZN(new_n244));
  AOI21_X1  g0044(.A(G1), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(new_n247), .A3(G274), .ZN(new_n248));
  INV_X1    g0048(.A(G226), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n248), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(G222), .B1(new_n261), .B2(G77), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n256), .B2(new_n257), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT66), .B(G223), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n247), .A2(KEYINPUT67), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n215), .B2(new_n246), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n253), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G190), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(new_n272), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  INV_X1    g0077(.A(G20), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n277), .A2(new_n278), .A3(G1), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n214), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n250), .B2(G20), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n284), .B2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(new_n201), .B2(new_n278), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT8), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n295));
  OAI21_X1  g0095(.A(G58), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT70), .B(G58), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n278), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n289), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n283), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n285), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n276), .B1(KEYINPUT9), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n308), .B(new_n311), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n272), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G169), .B2(new_n272), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(new_n307), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n256), .A2(new_n278), .A3(new_n257), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n278), .A4(new_n257), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n290), .A2(new_n322), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G159), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n288), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n321), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT76), .B1(new_n259), .B2(new_n260), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n256), .A2(new_n335), .A3(new_n257), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(new_n278), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n324), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n322), .B1(new_n338), .B2(new_n326), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n332), .A2(new_n321), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n333), .B(new_n283), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n300), .A2(new_n279), .ZN(new_n342));
  INV_X1    g0142(.A(new_n284), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n300), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  OAI211_X1 g0147(.A(G223), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n348));
  OAI211_X1 g0148(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n271), .ZN(new_n352));
  INV_X1    g0152(.A(new_n252), .ZN(new_n353));
  INV_X1    g0153(.A(G274), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n215), .B2(new_n246), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(G232), .B1(new_n355), .B2(new_n245), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n347), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G232), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n248), .B1(new_n359), .B2(new_n252), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n271), .B2(new_n351), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n346), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT18), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n341), .A2(new_n345), .B1(new_n358), .B2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n352), .A2(new_n356), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n361), .B2(G200), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n341), .A2(new_n345), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n341), .A2(new_n371), .A3(KEYINPUT17), .A4(new_n345), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n365), .A2(new_n368), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n303), .A2(G77), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n322), .A2(G20), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G50), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n288), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n283), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT11), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT11), .B(new_n283), .C1(new_n383), .C2(new_n384), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n279), .A2(KEYINPUT75), .A3(new_n322), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT12), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n280), .B2(G68), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n392), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(G68), .B2(new_n284), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n258), .A2(G226), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G97), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT3), .B(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(G232), .A3(G1698), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n271), .ZN(new_n402));
  INV_X1    g0202(.A(new_n248), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(G238), .B2(new_n353), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(G169), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(G179), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n410), .B1(new_n409), .B2(G169), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n396), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n388), .A2(new_n395), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(G190), .A3(new_n408), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n409), .A2(G200), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n387), .A4(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n353), .A2(G244), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n264), .A2(G238), .B1(new_n261), .B2(G107), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n399), .A2(G232), .A3(new_n263), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI211_X1 g0223(.A(new_n403), .B(new_n420), .C1(new_n271), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n316), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n284), .A2(G77), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G77), .B2(new_n280), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT8), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G58), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n291), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n301), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n434), .B2(new_n283), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n425), .B(new_n436), .C1(G169), .C2(new_n424), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n424), .A2(G190), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n435), .C1(new_n275), .C2(new_n424), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n377), .A2(new_n415), .A3(new_n419), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n320), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n325), .A2(new_n326), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(G107), .B1(G77), .B2(new_n287), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT77), .ZN(new_n446));
  AND2_X1   g0246(.A1(G97), .A2(G107), .ZN(new_n447));
  NOR2_X1   g0247(.A1(G97), .A2(G107), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT78), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G97), .A2(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n206), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT6), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n283), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  OAI211_X1 g0259(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n460));
  OAI211_X1 g0260(.A(G244), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT4), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT4), .B1(new_n258), .B2(G244), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n271), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n247), .A2(G274), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n244), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n468), .A2(new_n469), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n467), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(G257), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n280), .A2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n250), .A2(G33), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n280), .A2(new_n305), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(G97), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n465), .A2(new_n475), .A3(G190), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n458), .A2(new_n477), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n465), .A2(G179), .A3(new_n475), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n347), .B1(new_n465), .B2(new_n475), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n305), .B1(new_n444), .B2(new_n456), .ZN(new_n486));
  INV_X1    g0286(.A(new_n481), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT79), .B1(new_n244), .B2(G1), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT79), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n250), .A3(G45), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n247), .A2(new_n490), .A3(new_n492), .A4(G250), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n247), .A2(G274), .A3(new_n467), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT80), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n499));
  OAI211_X1 g0299(.A(G238), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n496), .A2(new_n498), .B1(new_n271), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G190), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n271), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n497), .B1(new_n493), .B2(new_n494), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n399), .A2(new_n278), .A3(G68), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n278), .B1(new_n398), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(G87), .B2(new_n206), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n301), .B2(new_n204), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n283), .B1(new_n279), .B2(new_n433), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n480), .A2(G87), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n504), .A2(new_n509), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n433), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n480), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n508), .A2(new_n347), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n503), .A2(new_n316), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n470), .A2(G264), .A3(new_n247), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT84), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n399), .A2(new_n528), .A3(G257), .A4(G1698), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n525), .B1(new_n532), .B2(new_n271), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n473), .A2(new_n355), .A3(new_n467), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n316), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n530), .B(new_n531), .C1(new_n526), .C2(KEYINPUT84), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n528), .B1(new_n264), .B2(G257), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n271), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n525), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n347), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n278), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n399), .A2(new_n544), .A3(new_n278), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n501), .A2(G20), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n278), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT24), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n305), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT25), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n280), .B2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n480), .A2(G107), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n535), .B(new_n541), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n546), .B2(new_n551), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n283), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n540), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n533), .A2(G190), .A3(new_n534), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n560), .A4(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n489), .A2(new_n524), .A3(new_n562), .A4(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n263), .A2(G264), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G257), .A2(G1698), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n570), .A2(new_n571), .B1(new_n259), .B2(new_n260), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n247), .A2(KEYINPUT67), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n215), .A2(new_n269), .A3(new_n246), .ZN(new_n574));
  INV_X1    g0374(.A(G303), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n256), .A2(new_n575), .A3(new_n257), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(new_n534), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n470), .A2(G270), .A3(new_n247), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT81), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n470), .A2(new_n581), .A3(G270), .A4(new_n247), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n578), .B2(new_n583), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n282), .A2(new_n214), .B1(G20), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n459), .B(new_n278), .C1(G33), .C2(new_n204), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n588), .B2(new_n589), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n279), .A2(new_n587), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n280), .A2(new_n305), .A3(new_n479), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(new_n587), .ZN(new_n596));
  OAI21_X1  g0396(.A(G169), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n585), .A2(new_n586), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT21), .B1(new_n598), .B2(KEYINPUT83), .ZN(new_n599));
  OAI21_X1  g0399(.A(G190), .B1(new_n585), .B2(new_n586), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n591), .A2(new_n592), .ZN(new_n601));
  INV_X1    g0401(.A(new_n594), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n480), .B2(G116), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n578), .A2(new_n583), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT82), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n600), .B(new_n605), .C1(new_n609), .C2(new_n275), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n347), .B1(new_n601), .B2(new_n603), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n578), .A2(new_n583), .A3(G179), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n605), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n599), .A2(new_n610), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n569), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n442), .A2(new_n620), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n365), .A2(new_n368), .ZN(new_n622));
  INV_X1    g0422(.A(new_n419), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n415), .B1(new_n623), .B2(new_n437), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n374), .A2(new_n375), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n314), .A2(new_n315), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n319), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n599), .A2(new_n615), .A3(new_n618), .A4(new_n562), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n483), .A2(new_n488), .A3(new_n523), .A4(new_n518), .ZN(new_n632));
  INV_X1    g0432(.A(new_n568), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(new_n485), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n465), .A2(new_n475), .A3(G179), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT85), .B1(new_n484), .B2(new_n485), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n458), .A2(new_n481), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n518), .A2(new_n523), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n488), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n524), .A2(new_n646), .A3(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n635), .A2(new_n648), .A3(new_n523), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n442), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n630), .A2(new_n650), .ZN(G369));
  INV_X1    g0451(.A(G330), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n614), .B1(new_n612), .B2(new_n613), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n617), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n250), .A2(new_n278), .A3(G13), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT86), .B(G343), .Z(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n605), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n619), .A2(new_n665), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n652), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n562), .A2(new_n664), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT87), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n562), .A2(KEYINPUT87), .A3(new_n664), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n562), .A2(new_n568), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n664), .B1(new_n565), .B2(new_n560), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n671), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n655), .A2(new_n663), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n562), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n664), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n209), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n212), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(new_n523), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n631), .B2(new_n634), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n486), .A2(new_n487), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n637), .A2(new_n639), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(KEYINPUT85), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n524), .A2(new_n694), .A3(KEYINPUT26), .A4(new_n640), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n636), .B1(new_n644), .B2(new_n488), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n663), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n663), .B1(new_n691), .B2(new_n648), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  INV_X1    g0502(.A(new_n476), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n577), .A2(new_n534), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n580), .B2(new_n582), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT89), .B1(new_n705), .B2(G179), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n578), .A2(new_n583), .A3(KEYINPUT89), .A4(G179), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n703), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n538), .A2(new_n539), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT88), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n508), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT88), .B1(new_n503), .B2(new_n533), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n702), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n616), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n476), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n711), .B1(new_n710), .B2(new_n508), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n503), .A2(new_n533), .A3(KEYINPUT88), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n540), .A2(new_n476), .A3(new_n316), .A4(new_n508), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n609), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n715), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n663), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n632), .A2(new_n673), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n655), .A2(new_n610), .A3(new_n730), .A4(new_n664), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n701), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n689), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(new_n277), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n250), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n684), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n668), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n666), .A2(new_n667), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n652), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n214), .B1(G20), .B2(new_n347), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n278), .A2(new_n316), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n369), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n278), .A2(new_n369), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n316), .A2(G200), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n754), .A2(new_n382), .B1(new_n290), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n278), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n759), .B1(G77), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT92), .Z(new_n768));
  NOR2_X1   g0568(.A1(new_n275), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G87), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n399), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(new_n760), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n205), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(KEYINPUT93), .B2(new_n772), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n278), .B1(new_n780), .B2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n204), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n760), .A2(new_n780), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G159), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(new_n785), .B2(KEYINPUT32), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(KEYINPUT32), .B2(new_n785), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT95), .ZN(new_n788));
  INV_X1    g0588(.A(new_n752), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n369), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n752), .A2(KEYINPUT95), .A3(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n787), .B1(new_n793), .B2(G68), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n768), .A2(new_n773), .A3(new_n779), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n770), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G303), .A2(new_n798), .B1(new_n784), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n261), .C1(new_n800), .C2(new_n758), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n797), .B(new_n801), .C1(G326), .C2(new_n753), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n777), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G283), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n766), .A2(G311), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n804), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n750), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n747), .A2(new_n749), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n334), .A2(new_n336), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n683), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n213), .A2(new_n244), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n238), .C2(new_n244), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n683), .A2(new_n261), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G355), .B1(new_n587), .B2(new_n683), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT90), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n810), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  INV_X1    g0620(.A(new_n740), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n809), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n748), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n744), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n749), .A2(new_n745), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G107), .A2(new_n798), .B1(new_n784), .B2(G311), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n261), .C1(new_n796), .C2(new_n758), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n782), .B(new_n829), .C1(G303), .C2(new_n753), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n777), .A2(new_n771), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G116), .B2(new_n766), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n830), .B(new_n832), .C1(new_n833), .C2(new_n792), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT96), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n766), .A2(G159), .B1(G143), .B2(new_n757), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n792), .A2(new_n286), .B1(new_n837), .B2(new_n754), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT97), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n777), .A2(new_n322), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G50), .A2(new_n798), .B1(new_n784), .B2(G132), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n811), .C1(new_n290), .C2(new_n781), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(new_n842), .C2(new_n843), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n835), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n740), .B1(G77), .B2(new_n827), .C1(new_n849), .C2(new_n750), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT98), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n437), .A2(new_n663), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n439), .B1(new_n435), .B2(new_n664), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n437), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n852), .B(new_n853), .C1(new_n745), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n440), .A2(new_n664), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n691), .B2(new_n648), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n700), .B2(new_n856), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n734), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n734), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n863), .A2(new_n864), .A3(new_n740), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n858), .A2(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n737), .A2(new_n250), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  INV_X1    g0668(.A(new_n859), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n854), .B1(new_n649), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n396), .A2(new_n663), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n415), .A2(new_n419), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n396), .B(new_n663), .C1(new_n413), .C2(new_n414), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n868), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT101), .B(new_n874), .C1(new_n860), .C2(new_n854), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n332), .A2(new_n321), .ZN(new_n878));
  INV_X1    g0678(.A(new_n326), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n337), .B2(new_n324), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(new_n322), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n283), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n321), .B1(new_n339), .B2(new_n332), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n882), .A2(new_n883), .B1(new_n342), .B2(new_n344), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n661), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n376), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT102), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n352), .A2(G179), .A3(new_n356), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n888), .A2(new_n357), .A3(new_n660), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n283), .A3(new_n881), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n345), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n341), .A2(new_n345), .A3(new_n371), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n887), .B(KEYINPUT37), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n346), .A2(new_n660), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n364), .A2(new_n894), .A3(new_n895), .A4(new_n372), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n372), .B1(new_n884), .B2(new_n889), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n887), .B1(new_n898), .B2(KEYINPUT37), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n886), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n886), .B(KEYINPUT38), .C1(new_n897), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n876), .A2(new_n877), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  INV_X1    g0706(.A(new_n903), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n892), .A2(new_n366), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT104), .A3(new_n895), .A4(new_n894), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n364), .A2(new_n894), .A3(new_n372), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n376), .A2(new_n346), .A3(new_n660), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n906), .B1(new_n907), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n396), .B(new_n664), .C1(new_n413), .C2(new_n414), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT103), .Z(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n622), .A2(new_n661), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n905), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n905), .A2(new_n922), .A3(KEYINPUT105), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n699), .B(new_n442), .C1(KEYINPUT29), .C2(new_n700), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n630), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n928), .B(new_n930), .Z(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n732), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n726), .A2(KEYINPUT106), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n620), .A2(new_n664), .B1(new_n727), .B2(new_n728), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n914), .A2(new_n915), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n901), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n903), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n874), .A2(new_n856), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n941), .B1(new_n935), .B2(new_n936), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n943), .A2(KEYINPUT40), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n937), .A2(new_n442), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n652), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n867), .B1(new_n931), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n931), .B2(new_n950), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n214), .A2(new_n278), .A3(new_n587), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT99), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(KEYINPUT35), .C2(new_n455), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT36), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT36), .ZN(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n290), .B2(new_n322), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n961), .A2(new_n212), .B1(G50), .B2(new_n322), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n277), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT100), .Z(new_n964));
  NAND4_X1  g0764(.A1(new_n952), .A2(new_n959), .A3(new_n960), .A4(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n489), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n692), .A2(new_n664), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(new_n643), .B2(new_n664), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT108), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n488), .B1(new_n970), .B2(new_n562), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n664), .ZN(new_n972));
  INV_X1    g0772(.A(new_n678), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n968), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT42), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n976), .A3(new_n968), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n516), .A2(new_n517), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n663), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n523), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n524), .A2(new_n980), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n978), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n676), .A2(new_n970), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n975), .A2(new_n977), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n994), .A2(new_n989), .A3(new_n988), .A4(new_n972), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n993), .B1(new_n992), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n684), .B(KEYINPUT41), .Z(new_n999));
  OAI211_X1 g0799(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n681), .C2(new_n968), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n678), .A2(new_n680), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n968), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n678), .A2(new_n680), .A3(new_n968), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT45), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n668), .B(new_n675), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1007), .B(KEYINPUT45), .Z(new_n1010));
  NAND4_X1  g0810(.A1(new_n1010), .A2(new_n676), .A3(new_n1000), .A4(new_n1005), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n675), .A2(new_n677), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n668), .A3(new_n678), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n742), .A2(new_n652), .B1(new_n973), .B2(new_n1012), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n735), .A2(KEYINPUT110), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n701), .A2(new_n734), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1009), .A2(new_n1011), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n999), .B1(new_n1021), .B2(new_n735), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n998), .B1(new_n1022), .B2(new_n739), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n812), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n234), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n810), .B1(new_n209), .B2(new_n433), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n740), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n774), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1028), .A2(G97), .B1(new_n784), .B2(G317), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n575), .B2(new_n758), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n781), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n811), .B(new_n1030), .C1(G107), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n770), .B2(new_n587), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n798), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1035));
  INV_X1    g0835(.A(G311), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1035), .C1(new_n754), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n793), .B2(G294), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1032), .B(new_n1038), .C1(new_n833), .C2(new_n765), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n792), .A2(new_n331), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n781), .A2(new_n322), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n399), .B1(new_n783), .B2(new_n837), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G143), .C2(new_n753), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n770), .A2(new_n290), .B1(new_n774), .B2(new_n202), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G150), .B2(new_n757), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n382), .C2(new_n765), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT47), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1027), .B1(new_n1048), .B2(new_n749), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n747), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n987), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1023), .A2(new_n1051), .ZN(G387));
  NAND3_X1  g0852(.A1(new_n1015), .A2(new_n739), .A3(new_n1014), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G77), .A2(new_n798), .B1(new_n784), .B2(G150), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n811), .B(new_n1054), .C1(new_n777), .C2(new_n204), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n793), .A2(new_n300), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G50), .A2(new_n757), .B1(new_n1031), .B2(new_n519), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT113), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n766), .A2(G68), .B1(G159), .B2(new_n753), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n811), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1028), .A2(G116), .B1(new_n784), .B2(G326), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n770), .A2(new_n796), .B1(new_n781), .B2(new_n833), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n753), .A2(G322), .B1(G317), .B2(new_n757), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n765), .B2(new_n575), .C1(new_n792), .C2(new_n1036), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT114), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1062), .B(new_n1063), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1061), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n749), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n686), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n815), .A2(new_n1076), .B1(new_n205), .B2(new_n683), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT111), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n230), .A2(new_n244), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n431), .A2(new_n382), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT50), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n686), .B(new_n244), .C1(new_n322), .C2(new_n202), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n812), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n821), .B1(new_n1084), .B2(new_n810), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1075), .B(new_n1085), .C1(new_n675), .C2(new_n1050), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n684), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1053), .B(new_n1086), .C1(new_n1087), .C2(new_n1089), .ZN(G393));
  NAND3_X1  g0890(.A1(new_n1009), .A2(new_n1011), .A3(new_n739), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n970), .A2(new_n747), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n753), .A2(G317), .B1(G311), .B2(new_n757), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n778), .B1(G294), .B2(new_n766), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n261), .B1(new_n783), .B2(new_n800), .C1(new_n833), .C2(new_n770), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G116), .B2(new_n1031), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(new_n575), .C2(new_n792), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n831), .B1(new_n431), .B2(new_n766), .ZN(new_n1099));
  INV_X1    g0899(.A(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n770), .A2(new_n322), .B1(new_n783), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n1062), .C1(G77), .C2(new_n1031), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1099), .B(new_n1102), .C1(new_n382), .C2(new_n792), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n753), .A2(G150), .B1(G159), .B2(new_n757), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT51), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1094), .A2(new_n1098), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT115), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n749), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n810), .B1(new_n204), .B2(new_n209), .C1(new_n1024), .C2(new_n241), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1092), .A2(new_n740), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1021), .A2(new_n684), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1011), .A2(new_n1009), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1091), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(G390));
  AOI21_X1  g0913(.A(new_n652), .B1(new_n935), .B2(new_n936), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n442), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n630), .A3(new_n929), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n937), .A2(G330), .A3(new_n942), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n718), .A2(new_n721), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n724), .B1(new_n1118), .B2(new_n702), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n664), .B1(new_n1119), .B2(new_n722), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n731), .B1(KEYINPUT31), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n732), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n856), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n875), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n870), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n937), .A2(G330), .A3(new_n856), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n875), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n733), .A2(G330), .A3(new_n856), .A4(new_n874), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n855), .A2(new_n437), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n854), .B1(new_n698), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1116), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1117), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n874), .B1(new_n860), .B2(new_n854), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n917), .A2(new_n921), .B1(new_n1138), .B2(new_n919), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n635), .A2(new_n697), .A3(new_n523), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n664), .A3(new_n1131), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n854), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n875), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n919), .B1(new_n907), .B2(new_n916), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1137), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n919), .B1(new_n870), .B2(new_n875), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT39), .B1(new_n939), .B2(new_n903), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n919), .B(new_n940), .C1(new_n1132), .C2(new_n875), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n1130), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1136), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1114), .A2(new_n942), .B1(new_n1123), .B2(new_n875), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n874), .B1(new_n1114), .B2(new_n856), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1155), .A2(new_n870), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1116), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n1152), .A3(new_n1146), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n684), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1153), .A2(new_n738), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n745), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n740), .B1(new_n300), .B2(new_n827), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1028), .A2(G50), .B1(new_n784), .B2(G125), .ZN(new_n1165));
  INV_X1    g0965(.A(G132), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n399), .C1(new_n1166), .C2(new_n758), .ZN(new_n1167));
  INV_X1    g0967(.A(G128), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n754), .A2(new_n1168), .B1(new_n781), .B2(new_n331), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n798), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT53), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n770), .B2(new_n286), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n766), .A2(new_n1172), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1170), .B(new_n1176), .C1(new_n837), .C2(new_n792), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n261), .B1(new_n770), .B2(new_n771), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n754), .A2(new_n833), .B1(new_n781), .B2(new_n202), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G116), .C2(new_n757), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n204), .B2(new_n765), .C1(new_n205), .C2(new_n792), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n845), .B1(G294), .B2(new_n784), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT116), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1164), .B1(new_n1184), .B2(new_n749), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1162), .B1(new_n1163), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1161), .A2(new_n1186), .ZN(G378));
  NOR2_X1   g0987(.A1(new_n307), .A2(new_n661), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n320), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n320), .A2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n946), .B2(new_n652), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n944), .A2(new_n945), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT40), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n944), .B2(new_n940), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1198), .B(G330), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1197), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n928), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1197), .A2(new_n926), .A3(new_n1202), .A4(new_n927), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n739), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n740), .B1(G50), .B2(new_n827), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n774), .A2(new_n290), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G283), .B2(new_n784), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n202), .B2(new_n770), .C1(new_n205), .C2(new_n758), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1041), .B(new_n1210), .C1(G116), .C2(new_n753), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1062), .A2(new_n243), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n766), .B2(new_n519), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n204), .C2(new_n792), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G50), .B1(new_n255), .B2(new_n243), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1214), .A2(new_n1215), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n781), .A2(new_n286), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n758), .A2(new_n1168), .B1(new_n770), .B2(new_n1171), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G125), .C2(new_n753), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n1166), .B2(new_n792), .C1(new_n837), .C2(new_n765), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  OR2_X1    g1023(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n784), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(new_n255), .A3(new_n243), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1223), .B(new_n1227), .C1(new_n331), .C2(new_n774), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1217), .B1(new_n1215), .B2(new_n1214), .C1(new_n1222), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1207), .B1(new_n1229), .B2(new_n749), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1198), .B2(new_n746), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1206), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1126), .A2(new_n1125), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1234));
  OAI211_X1 g1034(.A(KEYINPUT118), .B(new_n1159), .C1(new_n1153), .C2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT118), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n684), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1159), .B1(new_n1153), .B2(new_n1234), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT118), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1235), .ZN(new_n1244));
  AND4_X1   g1044(.A1(new_n926), .A2(new_n1197), .A3(new_n927), .A4(new_n1202), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1197), .A2(new_n1202), .B1(new_n926), .B2(new_n927), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1233), .B1(new_n1240), .B2(new_n1248), .ZN(G375));
  NAND3_X1  g1049(.A1(new_n1127), .A2(new_n1134), .A3(new_n1116), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n999), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1136), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(KEYINPUT119), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(KEYINPUT119), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n738), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n875), .A2(new_n745), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n740), .B1(G68), .B2(new_n827), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT120), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n793), .A2(new_n1172), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n811), .B1(new_n382), .B2(new_n781), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G132), .B2(new_n753), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n766), .A2(G150), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n770), .A2(new_n331), .B1(new_n783), .B2(new_n1168), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1208), .B(new_n1264), .C1(G137), .C2(new_n757), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G107), .A2(new_n766), .B1(new_n805), .B2(G77), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n261), .B1(new_n783), .B2(new_n575), .C1(new_n204), .C2(new_n770), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G294), .B2(new_n753), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1267), .B(new_n1269), .C1(new_n587), .C2(new_n792), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G283), .A2(new_n757), .B1(new_n1031), .B2(new_n519), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT121), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1266), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1259), .B1(new_n1273), .B2(new_n749), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1257), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1255), .B1(new_n1256), .B2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(KEYINPUT122), .B(new_n1275), .C1(new_n1234), .C2(new_n738), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1253), .A2(new_n1254), .A3(new_n1279), .ZN(G381));
  NOR3_X1   g1080(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1023), .A4(new_n1051), .ZN(new_n1283));
  OR3_X1    g1083(.A1(new_n1283), .A2(G378), .A3(G381), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G375), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT123), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1284), .A2(KEYINPUT123), .A3(G375), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G407));
  INV_X1    g1089(.A(G378), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n662), .A2(G213), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT124), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT125), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  OAI221_X1 g1094(.A(G213), .B1(G375), .B2(new_n1294), .C1(new_n1287), .C2(new_n1288), .ZN(G409));
  NAND3_X1  g1095(.A1(new_n1023), .A2(G390), .A3(new_n1051), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n824), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(new_n1282), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(KEYINPUT127), .A3(new_n1296), .A4(new_n1299), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G378), .B(new_n1233), .C1(new_n1240), .C2(new_n1248), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1244), .A2(new_n1247), .A3(new_n1251), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1290), .B1(new_n1307), .B2(new_n1232), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1292), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1250), .B1(new_n1135), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1116), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n684), .A3(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1314), .A2(new_n1279), .A3(G384), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1314), .B2(new_n1279), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1309), .A2(new_n1310), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1293), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1279), .ZN(new_n1321));
  INV_X1    g1121(.A(G384), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1314), .A2(new_n1279), .A3(G384), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(new_n1319), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1318), .A2(new_n1319), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(G2897), .A3(new_n1293), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1292), .A2(G2897), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT126), .B1(new_n1317), .B2(new_n1330), .ZN(new_n1331));
  AND4_X1   g1131(.A1(KEYINPUT126), .A2(new_n1323), .A3(new_n1324), .A4(new_n1330), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1329), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1328), .B1(new_n1333), .B2(new_n1320), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1305), .B1(new_n1327), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1305), .A2(KEYINPUT61), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1323), .A2(new_n1324), .A3(new_n1330), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT126), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1338), .B(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1337), .A2(new_n1340), .A3(new_n1329), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1318), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1336), .A2(new_n1341), .A3(new_n1343), .A4(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1335), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1290), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1306), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1317), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1347), .A2(new_n1325), .A3(new_n1306), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1305), .ZN(G402));
endmodule


