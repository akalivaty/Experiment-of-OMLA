//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT22), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G110), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G119), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n193), .A2(KEYINPUT76), .A3(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT76), .B1(new_n193), .B2(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n192), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT75), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n195), .B1(new_n210), .B2(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n201), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n198), .A2(new_n192), .A3(new_n200), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n211), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n191), .B1(new_n220), .B2(KEYINPUT77), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n213), .B2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n222), .B(new_n191), .C1(new_n213), .C2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT74), .B(G902), .Z(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n187), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g044(.A(KEYINPUT25), .B(new_n227), .C1(new_n224), .C2(new_n225), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n228), .B2(G234), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(G902), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT78), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT32), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n246), .A3(new_n249), .A4(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(new_n206), .B2(G143), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n254), .A3(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n199), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n206), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(G146), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n263), .B1(KEYINPUT0), .B2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n199), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n259), .A2(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n248), .A2(KEYINPUT67), .A3(new_n250), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT66), .A2(G119), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT66), .A2(G119), .ZN(new_n270));
  OAI21_X1  g084(.A(G116), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G119), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT2), .B(G113), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n256), .A2(new_n258), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n199), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n262), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  OAI21_X1  g097(.A(G128), .B1(new_n255), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n262), .A2(new_n263), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n244), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n242), .A2(G137), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n250), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n268), .A2(new_n279), .A3(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT26), .B(G101), .Z(new_n293));
  NOR2_X1   g107(.A1(G237), .A2(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G210), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n268), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n266), .A2(new_n251), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n279), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n292), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n300), .A2(KEYINPUT31), .A3(new_n307), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n292), .B(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n306), .A2(new_n303), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n298), .B(KEYINPUT70), .Z(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G472), .A2(G902), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT71), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n240), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n312), .A2(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n325), .A2(KEYINPUT32), .A3(new_n322), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n325), .A2(new_n322), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n324), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT72), .A3(new_n240), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n317), .A2(new_n318), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n307), .A2(new_n292), .ZN(new_n334));
  INV_X1    g148(.A(new_n298), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n268), .A2(new_n291), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n306), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n315), .A2(KEYINPUT29), .A3(new_n298), .A4(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  OAI221_X1 g158(.A(new_n228), .B1(new_n333), .B2(new_n338), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G472), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n239), .B1(new_n332), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT9), .B(G234), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G221), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n352));
  INV_X1    g166(.A(G104), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n353), .B2(G107), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n355));
  INV_X1    g169(.A(G107), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G104), .ZN(new_n357));
  INV_X1    g171(.A(G101), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(G107), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n354), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n356), .A2(G104), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n353), .A2(G107), .ZN(new_n362));
  OAI21_X1  g176(.A(G101), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(new_n287), .A3(KEYINPUT10), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n372), .A3(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n266), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n280), .A2(new_n262), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n199), .A2(KEYINPUT79), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n281), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n360), .A2(new_n363), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n284), .B1(new_n259), .B2(new_n377), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(KEYINPUT80), .A3(new_n383), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n375), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n253), .A2(new_n267), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n382), .A2(KEYINPUT80), .A3(new_n383), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT80), .B1(new_n382), .B2(new_n383), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT82), .B1(new_n394), .B2(new_n375), .ZN(new_n395));
  AND4_X1   g209(.A1(KEYINPUT82), .A2(new_n375), .A3(new_n386), .A4(new_n387), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n388), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n375), .A2(new_n386), .A3(KEYINPUT82), .A4(new_n387), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT83), .A3(new_n390), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n391), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n188), .A2(G227), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  OAI21_X1  g222(.A(new_n352), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n391), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT83), .B1(new_n403), .B2(new_n390), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n398), .B(new_n389), .C1(new_n401), .C2(new_n402), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT84), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n391), .A2(new_n414), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n382), .B1(new_n287), .B2(new_n380), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT12), .B1(new_n418), .B2(new_n390), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n418), .A2(new_n251), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(KEYINPUT12), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(new_n415), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n228), .ZN(new_n426));
  INV_X1    g240(.A(G902), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n417), .B1(new_n399), .B2(new_n404), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n414), .B1(new_n421), .B2(new_n391), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n432), .B2(G469), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n351), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n287), .A2(G125), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n266), .A2(new_n202), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G224), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n440), .A2(new_n445), .A3(new_n442), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  XOR2_X1   g264(.A(G110), .B(G122), .Z(new_n451));
  OAI211_X1 g265(.A(new_n373), .B(new_n371), .C1(new_n277), .C2(new_n278), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n271), .A2(KEYINPUT5), .A3(new_n273), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n453), .B(G113), .C1(KEYINPUT5), .C2(new_n271), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n274), .A2(new_n276), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n365), .A4(new_n367), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n452), .B2(new_n456), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n456), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n451), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n450), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n451), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n458), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT6), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n449), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT87), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n454), .A2(new_n455), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n364), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n451), .B(KEYINPUT8), .Z(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n438), .A2(KEYINPUT7), .A3(new_n446), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n439), .B1(new_n479), .B2(new_n445), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n464), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n427), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n470), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n473), .B1(new_n470), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n435), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(G475), .A2(G902), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT92), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n204), .B(KEYINPUT89), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n215), .B1(new_n490), .B2(new_n206), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n294), .A2(G214), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT88), .A3(G143), .ZN(new_n493));
  OR2_X1    g307(.A1(KEYINPUT88), .A2(G143), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT88), .A2(G143), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(G214), .A3(new_n294), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n496), .A3(G131), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n498), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n249), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n491), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT19), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n204), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n206), .B(new_n505), .C1(new_n490), .C2(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT90), .A3(new_n214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n497), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT90), .B1(new_n506), .B2(new_n214), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n353), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n207), .B(new_n517), .C1(new_n508), .C2(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n503), .A3(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT91), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n518), .A2(new_n503), .A3(new_n521), .A4(new_n513), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT20), .B(new_n489), .C1(new_n515), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n511), .A2(new_n514), .B1(new_n520), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n488), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n518), .B2(new_n503), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n520), .B2(new_n522), .ZN(new_n529));
  OAI21_X1  g343(.A(G475), .B1(new_n529), .B2(G902), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n349), .A2(new_n233), .A3(G953), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n254), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n199), .A2(G143), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G128), .B(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n539), .A3(new_n242), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(G134), .C1(KEYINPUT13), .C2(new_n533), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n272), .A2(G122), .ZN(new_n543));
  INV_X1    g357(.A(G122), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G116), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT93), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT93), .ZN(new_n548));
  AOI21_X1  g362(.A(G107), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n548), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n550), .A2(new_n356), .A3(new_n546), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n540), .B(new_n542), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n356), .B1(new_n550), .B2(new_n546), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT14), .B1(new_n544), .B2(G116), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT95), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n543), .A2(new_n557), .A3(KEYINPUT14), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n544), .A2(KEYINPUT14), .A3(G116), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n559), .A4(new_n545), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G107), .ZN(new_n561));
  INV_X1    g375(.A(new_n540), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n242), .B1(new_n537), .B2(new_n539), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n554), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n561), .A2(new_n554), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n537), .A2(new_n539), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G134), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n540), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(KEYINPUT96), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n553), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n532), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n564), .A2(new_n565), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT96), .B1(new_n567), .B2(new_n570), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n552), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(KEYINPUT97), .A3(new_n532), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n228), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n581), .A2(new_n583), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n531), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G952), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G953), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(G234), .B2(G237), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n188), .B(new_n228), .C1(G234), .C2(G237), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT21), .B(G898), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n486), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n347), .A2(new_n434), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(new_n239), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n325), .B2(new_n227), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n330), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n434), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n470), .A2(new_n483), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n471), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n470), .A2(new_n472), .A3(new_n483), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(new_n435), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n579), .A2(new_n607), .A3(new_n580), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n532), .B1(new_n577), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n532), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n572), .A2(KEYINPUT98), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n608), .A2(G478), .A3(new_n613), .A4(new_n228), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n581), .A2(new_n582), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n594), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n602), .A2(new_n606), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  AOI21_X1  g437(.A(new_n618), .B1(new_n585), .B2(new_n584), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n594), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n602), .A2(new_n606), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT35), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n356), .ZN(G9));
  NOR2_X1   g443(.A1(new_n586), .A2(new_n594), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n191), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n220), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n237), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n235), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n435), .ZN(new_n636));
  INV_X1    g450(.A(new_n473), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n603), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n470), .A2(new_n473), .A3(new_n483), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n630), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n434), .A2(new_n601), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n192), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AOI22_X1  g459(.A1(new_n329), .A2(new_n331), .B1(G472), .B2(new_n345), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n229), .A2(new_n231), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n647), .A2(new_n234), .B1(new_n237), .B2(new_n633), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n585), .A2(new_n584), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n590), .B1(new_n591), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n650), .A2(new_n531), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n624), .A2(KEYINPUT100), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n649), .A2(new_n434), .A3(new_n606), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  NAND2_X1  g475(.A1(new_n638), .A2(new_n639), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT38), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT38), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n618), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n318), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n292), .B2(new_n340), .ZN(new_n671));
  INV_X1    g485(.A(new_n310), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n427), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n332), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n636), .A3(new_n635), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n652), .B(KEYINPUT39), .Z(new_n677));
  AND2_X1   g491(.A1(new_n434), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n669), .B(new_n676), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  AOI21_X1  g496(.A(new_n531), .B1(new_n615), .B2(new_n614), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n653), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n649), .A2(new_n434), .A3(new_n606), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AND3_X1   g501(.A1(new_n424), .A2(new_n425), .A3(new_n228), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n425), .B1(new_n424), .B2(new_n228), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n604), .A2(new_n435), .A3(new_n605), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n351), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n347), .A3(new_n620), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n347), .A3(new_n626), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND3_X1  g510(.A1(new_n691), .A2(new_n630), .A3(new_n649), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NOR3_X1   g512(.A1(new_n688), .A2(new_n689), .A3(new_n351), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n315), .A2(new_n340), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n314), .B1(new_n700), .B2(new_n670), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n323), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n599), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n239), .A2(new_n594), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n668), .A2(new_n690), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n699), .A2(KEYINPUT102), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n424), .A2(new_n228), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n350), .A3(new_n426), .A4(new_n705), .ZN(new_n710));
  INV_X1    g524(.A(new_n704), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n544), .ZN(G24));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n648), .B2(new_n703), .ZN(new_n716));
  INV_X1    g530(.A(new_n703), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n635), .A2(new_n717), .A3(KEYINPUT103), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n684), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n699), .A2(new_n719), .A3(new_n606), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND3_X1  g535(.A1(new_n320), .A2(new_n240), .A3(new_n323), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT32), .B1(new_n325), .B2(new_n322), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n239), .B1(new_n727), .B2(new_n346), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n662), .A2(new_n636), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n684), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(new_n434), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n347), .A2(new_n434), .A3(new_n729), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(KEYINPUT105), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND2_X1  g555(.A1(new_n658), .A2(KEYINPUT106), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n347), .A2(new_n742), .A3(new_n434), .A4(new_n729), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n658), .A2(KEYINPUT106), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  OAI21_X1  g560(.A(new_n416), .B1(new_n411), .B2(new_n412), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT45), .A3(new_n430), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n429), .B2(new_n431), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n747), .A2(new_n752), .A3(KEYINPUT45), .A4(new_n430), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n749), .A2(G469), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n428), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n755), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n426), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n350), .A3(new_n677), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n616), .A2(new_n531), .ZN(new_n762));
  NAND2_X1  g576(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n600), .A3(new_n635), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n730), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n761), .B(new_n769), .C1(new_n768), .C2(new_n767), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  AND2_X1   g585(.A1(new_n646), .A2(new_n239), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n688), .B1(new_n756), .B2(new_n757), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n773), .B(new_n351), .C1(new_n774), .C2(new_n759), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n760), .B2(new_n350), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n731), .B(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT112), .B1(new_n775), .B2(new_n776), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n755), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n754), .B2(new_n755), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n688), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n773), .B1(new_n783), .B2(new_n351), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n350), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n688), .A2(new_n689), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT109), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n351), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n780), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n590), .A2(new_n766), .A3(new_n598), .A4(new_n717), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n729), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n699), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n665), .A2(new_n636), .A3(new_n666), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n798), .B2(new_n799), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n699), .A2(new_n729), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n716), .A2(new_n718), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n766), .A2(new_n590), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n675), .A2(new_n598), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n805), .A2(new_n590), .A3(new_n531), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n810), .B2(new_n616), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n792), .A2(new_n796), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(KEYINPUT113), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT51), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT115), .B1(new_n798), .B2(new_n690), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n794), .A2(new_n699), .A3(new_n817), .A4(new_n606), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n683), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n805), .A2(new_n590), .A3(new_n809), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n819), .B(new_n588), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n699), .A2(new_n807), .A3(new_n729), .A4(new_n728), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT48), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n815), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n821), .A2(new_n820), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n589), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n824), .A3(KEYINPUT116), .A4(new_n819), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(KEYINPUT114), .B(new_n808), .C1(new_n810), .C2(new_n616), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(KEYINPUT51), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n775), .A2(new_n776), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n795), .B1(new_n833), .B2(new_n791), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n811), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n835), .A3(new_n803), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n779), .B1(new_n814), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n831), .A2(new_n803), .A3(KEYINPUT51), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n834), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n837), .B1(new_n826), .B2(new_n829), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n797), .A2(new_n803), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n793), .B1(new_n792), .B2(new_n796), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n811), .ZN(new_n846));
  OAI211_X1 g660(.A(KEYINPUT117), .B(new_n843), .C1(new_n846), .C2(KEYINPUT51), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n692), .A2(new_n695), .A3(new_n697), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n713), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n683), .A2(new_n640), .A3(KEYINPUT110), .A4(new_n617), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n619), .B2(new_n486), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n640), .A2(new_n617), .A3(new_n624), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n434), .A2(new_n855), .A3(new_n598), .A4(new_n601), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n596), .A3(new_n642), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n856), .A2(new_n596), .A3(new_n642), .A4(KEYINPUT111), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n606), .A2(new_n650), .A3(new_n618), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n332), .B2(new_n674), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n434), .A3(new_n648), .A4(new_n653), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n720), .A2(new_n660), .A3(new_n686), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n646), .A2(new_n658), .A3(new_n648), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n351), .B(new_n690), .C1(new_n426), .C2(new_n433), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n691), .A2(new_n719), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n686), .A4(new_n864), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n850), .A2(new_n861), .A3(new_n866), .A4(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n586), .A2(new_n652), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n646), .A2(new_n648), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n434), .B(new_n729), .C1(new_n874), .C2(new_n719), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n744), .B2(new_n743), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n738), .B2(new_n739), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n848), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n692), .A2(new_n695), .A3(new_n697), .ZN(new_n881));
  INV_X1    g695(.A(new_n713), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n861), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n866), .A2(new_n871), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n876), .A2(new_n848), .A3(new_n736), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n879), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n866), .A2(new_n871), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n880), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n847), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n587), .A2(new_n188), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n789), .A2(new_n790), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT49), .Z(new_n898));
  INV_X1    g712(.A(new_n667), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n636), .A3(new_n762), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n350), .A3(new_n809), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(G75));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n879), .A2(new_n887), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n227), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n471), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT6), .B1(new_n468), .B2(new_n463), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n461), .A2(new_n450), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n449), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n188), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n903), .B(new_n911), .C1(new_n905), .C2(new_n471), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(G51));
  INV_X1    g731(.A(new_n754), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n904), .A2(new_n227), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n755), .A2(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n880), .B1(new_n879), .B2(new_n887), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n888), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n755), .A2(KEYINPUT57), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n424), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n914), .B1(new_n921), .B2(new_n926), .ZN(G54));
  NAND4_X1  g741(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .A4(new_n227), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(new_n526), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n526), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n914), .ZN(G60));
  AND2_X1   g745(.A1(new_n608), .A2(new_n613), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n932), .B(new_n935), .C1(new_n888), .C2(new_n923), .ZN(new_n936));
  INV_X1    g750(.A(new_n892), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n885), .A2(new_n877), .A3(new_n861), .A4(new_n850), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n938), .A2(new_n848), .B1(new_n890), .B2(new_n886), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n880), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n915), .B(new_n936), .C1(new_n941), .C2(new_n932), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(G63));
  INV_X1    g757(.A(new_n226), .ZN(new_n944));
  XOR2_X1   g758(.A(KEYINPUT119), .B(KEYINPUT60), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT120), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n939), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n904), .A2(new_n633), .A3(new_n948), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n951), .A3(new_n915), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(KEYINPUT121), .A3(new_n915), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT61), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n949), .B1(new_n879), .B2(new_n887), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n914), .B1(new_n955), .B2(new_n633), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n956), .B(new_n950), .C1(KEYINPUT121), .C2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n954), .A2(new_n958), .ZN(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n593), .B2(new_n444), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n884), .B2(G953), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n907), .B(new_n908), .C1(G898), .C2(new_n188), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n301), .A2(new_n305), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT122), .Z(new_n965));
  OAI21_X1  g779(.A(new_n505), .B1(new_n490), .B2(new_n504), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n820), .A2(new_n625), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n678), .A2(new_n347), .A3(new_n729), .A4(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n777), .A2(new_n770), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n869), .A2(KEYINPUT123), .A3(new_n686), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n720), .A2(new_n660), .A3(new_n686), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n681), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n972), .A2(new_n975), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .A3(new_n681), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n971), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n968), .B1(new_n981), .B2(G953), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n761), .A2(new_n705), .A3(new_n728), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n777), .A2(new_n770), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n987), .A2(new_n988), .A3(new_n740), .A4(new_n745), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n967), .B(new_n985), .C1(new_n989), .C2(G953), .ZN(new_n990));
  OAI211_X1 g804(.A(KEYINPUT124), .B(new_n968), .C1(new_n981), .C2(G953), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n984), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n984), .A2(new_n995), .A3(new_n990), .A4(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  XNOR2_X1  g811(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n981), .B2(new_n884), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n298), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n334), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1000), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n989), .B2(new_n883), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(new_n335), .A3(new_n292), .A4(new_n307), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n891), .A2(new_n879), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n336), .B(KEYINPUT127), .Z(new_n1011));
  OAI211_X1 g825(.A(new_n1010), .B(new_n1007), .C1(new_n672), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1009), .A2(new_n915), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1006), .A2(new_n1013), .ZN(G57));
endmodule


