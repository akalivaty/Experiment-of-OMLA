//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n206), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n209), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n224), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n211), .A2(new_n213), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n211), .A2(new_n213), .A3(new_n254), .A4(new_n251), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G68), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n211), .A2(new_n213), .A3(new_n251), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n264), .A2(new_n202), .B1(new_n216), .B2(G68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n216), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n262), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT11), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n254), .ZN(new_n272));
  INV_X1    g0072(.A(G68), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n269), .A2(new_n270), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n261), .A2(new_n271), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT73), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n211), .B2(new_n213), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  OAI211_X1 g0091(.A(G226), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT69), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n285), .A2(new_n294), .A3(G226), .A4(new_n289), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G1), .A3(G13), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G238), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AND2_X1   g0103(.A1(G1), .A2(G13), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n281), .B1(new_n297), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n308), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n286), .A2(new_n287), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n295), .B2(new_n293), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n280), .C1(new_n312), .C2(new_n284), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n279), .B1(new_n314), .B2(G169), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI211_X1 g0116(.A(KEYINPUT14), .B(new_n316), .C1(new_n309), .C2(new_n313), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n297), .A2(new_n308), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT71), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(KEYINPUT13), .C1(new_n297), .C2(new_n308), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n328), .A3(G179), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n278), .B1(new_n318), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n309), .B2(new_n313), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(new_n277), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n323), .A2(new_n321), .B1(new_n325), .B2(new_n327), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(G190), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n256), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G50), .A3(new_n260), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(new_n266), .B1(new_n340), .B2(new_n264), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G20), .B2(new_n203), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n338), .B1(G50), .B2(new_n254), .C1(new_n342), .C2(new_n252), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT9), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n285), .A2(G222), .A3(new_n289), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n285), .A2(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G223), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n347), .B1(new_n267), .B2(new_n285), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n283), .ZN(new_n351));
  INV_X1    g0151(.A(new_n307), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G226), .B2(new_n301), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n345), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n354), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(new_n331), .B1(new_n343), .B2(new_n344), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT10), .Z(new_n359));
  OAI21_X1  g0159(.A(new_n343), .B1(new_n356), .B2(G169), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n360), .A2(KEYINPUT67), .B1(new_n361), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(KEYINPUT67), .B2(new_n360), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n299), .A2(G232), .A3(new_n300), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n307), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G226), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G1698), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G223), .B2(G1698), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n290), .A2(new_n291), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n370), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n367), .B1(new_n283), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n361), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n283), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n301), .A2(G232), .B1(new_n305), .B2(new_n306), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n361), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n381));
  AOI21_X1  g0181(.A(G169), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n377), .B(KEYINPUT75), .C1(new_n381), .C2(new_n382), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n285), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n273), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n223), .A2(new_n273), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n201), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n263), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n387), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n371), .B2(new_n216), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n290), .A2(new_n291), .A3(new_n388), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n395), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n401), .A3(new_n262), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n339), .B1(new_n253), .B2(G20), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(new_n337), .B1(new_n272), .B2(new_n339), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n385), .A2(new_n386), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n378), .A2(new_n379), .A3(new_n346), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n375), .B2(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n410));
  OR2_X1    g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(KEYINPUT76), .B2(KEYINPUT17), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n406), .A2(KEYINPUT18), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n385), .A2(new_n414), .A3(new_n386), .A4(new_n405), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n285), .A2(G232), .A3(new_n289), .ZN(new_n418));
  INV_X1    g0218(.A(G107), .ZN(new_n419));
  INV_X1    g0219(.A(G238), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n418), .B1(new_n419), .B2(new_n285), .C1(new_n348), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n283), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n352), .B1(G244), .B2(new_n301), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n316), .ZN(new_n425));
  INV_X1    g0225(.A(new_n339), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n266), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n262), .B1(new_n267), .B2(new_n272), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n422), .A2(new_n361), .A3(new_n423), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n425), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n422), .A2(G190), .A3(new_n423), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(G200), .B2(new_n424), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n336), .A2(new_n365), .A3(new_n417), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT6), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n440), .A2(new_n225), .A3(G107), .ZN(new_n441));
  XNOR2_X1  g0241(.A(G97), .B(G107), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n443), .A2(new_n216), .B1(new_n267), .B2(new_n264), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n419), .B1(new_n389), .B2(new_n390), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n262), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n254), .A2(G97), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n256), .B1(new_n253), .B2(G33), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G97), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT5), .B(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n305), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n453), .A2(new_n452), .B1(new_n304), .B2(new_n298), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n456), .B2(new_n226), .ZN(new_n457));
  OAI211_X1 g0257(.A(G244), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n458), .A2(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n459), .ZN(new_n464));
  OAI211_X1 g0264(.A(G250), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n457), .B1(new_n468), .B2(new_n283), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n450), .B1(new_n469), .B2(G169), .ZN(new_n470));
  AOI211_X1 g0270(.A(G179), .B(new_n457), .C1(new_n468), .C2(new_n283), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n439), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G238), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n473));
  OAI211_X1 g0273(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n283), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n299), .A2(G274), .A3(new_n452), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n253), .A2(G45), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(G250), .C1(new_n282), .C2(new_n210), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(G169), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n477), .A2(new_n361), .A3(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT79), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n476), .B2(new_n283), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n361), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n483), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n216), .B1(new_n287), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n373), .A2(new_n225), .A3(new_n419), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n216), .B(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n266), .B2(new_n225), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT80), .A4(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n262), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n428), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n448), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n428), .A2(new_n272), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n486), .A2(new_n331), .ZN(new_n505));
  AOI211_X1 g0305(.A(new_n346), .B(new_n481), .C1(new_n283), .C2(new_n476), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n448), .A2(G87), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n500), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n489), .A2(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n454), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(G257), .B2(new_n455), .ZN(new_n512));
  INV_X1    g0312(.A(new_n464), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n466), .B(new_n465), .C1(new_n458), .C2(new_n459), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT77), .B1(new_n458), .B2(new_n459), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n516), .B2(new_n284), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n316), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n469), .A2(new_n361), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT78), .A4(new_n450), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n469), .A2(G190), .ZN(new_n521));
  INV_X1    g0321(.A(new_n450), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n331), .C2(new_n469), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n472), .A2(new_n510), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n216), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n285), .A2(new_n216), .A3(G87), .A4(new_n526), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n475), .A2(G20), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n216), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n419), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(new_n530), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n262), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n448), .A2(G107), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT25), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n254), .B2(G107), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n254), .A2(new_n542), .A3(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT83), .B(new_n542), .C1(new_n254), .C2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n226), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(G250), .B2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G294), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n553), .A2(new_n371), .B1(new_n372), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n283), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT84), .B1(new_n455), .B2(G264), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT5), .A2(G41), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT5), .A2(G41), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n452), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT84), .A3(G264), .A4(new_n299), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n454), .B(new_n556), .C1(new_n557), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(KEYINPUT85), .A3(G169), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(G264), .A3(new_n299), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n561), .B1(new_n283), .B2(new_n555), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G179), .A3(new_n454), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT85), .B1(new_n563), .B2(G169), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n551), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n530), .A2(new_n536), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n537), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n549), .B1(new_n575), .B2(new_n262), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n563), .A2(G190), .ZN(new_n577));
  AOI21_X1  g0377(.A(G200), .B1(new_n568), .B2(new_n454), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(G33), .B2(G283), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n372), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(G20), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n262), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n262), .A3(KEYINPUT20), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n583), .B2(new_n272), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n253), .A2(G33), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n255), .A2(G116), .A3(new_n258), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n285), .A2(new_n596), .A3(G257), .A4(new_n289), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n371), .A2(G303), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n283), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n560), .A2(G270), .A3(new_n299), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n602), .A2(new_n454), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(G190), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n603), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n593), .B(new_n604), .C1(new_n606), .C2(new_n331), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  INV_X1    g0408(.A(new_n591), .ZN(new_n609));
  INV_X1    g0409(.A(new_n588), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT20), .B1(new_n584), .B2(new_n262), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n610), .A2(new_n611), .B1(G116), .B2(new_n254), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n606), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n602), .A2(new_n454), .A3(G179), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n600), .B2(new_n283), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n592), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n316), .B1(new_n589), .B2(new_n591), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT21), .A3(new_n605), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n607), .A2(new_n614), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n580), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n438), .A2(new_n524), .A3(new_n621), .ZN(G372));
  AOI211_X1 g0422(.A(G179), .B(new_n481), .C1(new_n283), .C2(new_n476), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT86), .B1(new_n623), .B2(new_n483), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n484), .B(new_n625), .C1(G169), .C2(new_n486), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n504), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n500), .A2(new_n503), .A3(new_n508), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n506), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n505), .A2(KEYINPUT87), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n486), .B2(new_n331), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n627), .A2(new_n504), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n564), .A2(new_n569), .ZN(new_n636));
  INV_X1    g0436(.A(new_n571), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n576), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n614), .A2(new_n617), .A3(new_n619), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n579), .B(new_n635), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n472), .A2(new_n520), .A3(new_n523), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n628), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n470), .A2(new_n471), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n635), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n489), .A2(new_n504), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n507), .A2(new_n509), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n472), .B2(new_n520), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(KEYINPUT26), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n438), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n411), .A2(new_n412), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n334), .A2(G190), .ZN(new_n654));
  INV_X1    g0454(.A(new_n333), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n434), .ZN(new_n657));
  INV_X1    g0457(.A(new_n315), .ZN(new_n658));
  INV_X1    g0458(.A(new_n317), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n329), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n278), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n653), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n405), .A2(new_n383), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(new_n414), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n359), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n363), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n651), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n253), .A2(new_n216), .A3(G13), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  OAI21_X1  g0472(.A(G213), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n619), .A2(new_n617), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT21), .B1(new_n618), .B2(new_n605), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n639), .A2(KEYINPUT89), .A3(new_n675), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n572), .B(new_n579), .C1(new_n576), .C2(new_n675), .ZN(new_n682));
  INV_X1    g0482(.A(new_n675), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n638), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n680), .A2(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n638), .A2(new_n675), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT90), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n681), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n593), .A2(new_n675), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n620), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n639), .A2(new_n695), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(G330), .A3(new_n690), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n694), .A2(new_n700), .ZN(G399));
  NOR2_X1   g0501(.A1(new_n492), .A2(G116), .ZN(new_n702));
  INV_X1    g0502(.A(G41), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n207), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(G1), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n219), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n650), .A2(new_n708), .A3(new_n675), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n635), .A2(new_n643), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n472), .A2(new_n520), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n510), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n675), .B1(new_n642), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n621), .A2(new_n524), .A3(new_n675), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  INV_X1    g0521(.A(new_n615), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n568), .A2(new_n601), .A3(new_n486), .A4(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT91), .B(new_n721), .C1(new_n517), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n567), .A2(new_n561), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(new_n486), .A3(new_n556), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n469), .A2(new_n727), .A3(new_n616), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT91), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n486), .A2(G179), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n517), .A2(new_n563), .A3(new_n605), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n469), .A2(new_n727), .A3(KEYINPUT30), .A4(new_n616), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n725), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n720), .B1(new_n734), .B2(new_n675), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n721), .B1(new_n517), .B2(new_n723), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n732), .A3(new_n731), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n719), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT92), .B1(new_n718), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT92), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n709), .A2(new_n743), .A3(new_n717), .A4(new_n740), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n707), .B1(new_n745), .B2(G1), .ZN(G364));
  AND2_X1   g0546(.A1(new_n216), .A2(G13), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT93), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n704), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n750), .A2(new_n253), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n699), .B2(G330), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n699), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n285), .A2(new_n207), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n207), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n246), .A2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n371), .A2(new_n207), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n451), .B2(new_n220), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n215), .B1(G20), .B2(new_n316), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT94), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n752), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n216), .A2(new_n361), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n216), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n770), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G311), .A2(new_n772), .B1(new_n775), .B2(G329), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n769), .A2(new_n346), .A3(G200), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n371), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n346), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n216), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n781), .A2(new_n554), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n773), .A2(new_n346), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n779), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n785), .A2(new_n331), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT96), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(KEYINPUT96), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n792), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n285), .B1(new_n777), .B2(new_n273), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n775), .A2(G159), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n787), .A2(new_n223), .B1(new_n802), .B2(KEYINPUT32), .ZN(new_n803));
  INV_X1    g0603(.A(new_n782), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(G87), .C2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G77), .ZN(new_n810));
  INV_X1    g0610(.A(new_n797), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G50), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n789), .A2(new_n419), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n781), .A2(new_n225), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(KEYINPUT32), .C2(new_n802), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n805), .A2(new_n810), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n800), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n768), .B1(new_n817), .B2(new_n762), .ZN(new_n818));
  INV_X1    g0618(.A(new_n765), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n699), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n754), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n650), .A2(new_n675), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n675), .B1(new_n430), .B2(new_n431), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT100), .Z(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n437), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n425), .A2(new_n432), .A3(new_n433), .A4(new_n683), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT101), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n675), .B(new_n830), .C1(new_n642), .C2(new_n649), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n741), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n752), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(KEYINPUT102), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n832), .A2(new_n833), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n741), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT102), .B1(new_n834), .B2(new_n835), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n762), .A2(new_n763), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n752), .B1(new_n842), .B2(G77), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT98), .Z(new_n844));
  INV_X1    g0644(.A(new_n762), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n797), .A2(new_n783), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n789), .A2(new_n373), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n814), .A2(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n848), .B1(new_n419), .B2(new_n782), .C1(new_n554), .C2(new_n787), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n808), .A2(new_n583), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n371), .B1(new_n774), .B2(new_n851), .C1(new_n777), .C2(new_n790), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n846), .A2(new_n849), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n777), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G143), .A2(new_n786), .B1(new_n854), .B2(G150), .ZN(new_n855));
  INV_X1    g0655(.A(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(new_n808), .B2(new_n856), .C1(new_n797), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT34), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n285), .B1(new_n774), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n202), .A2(new_n782), .B1(new_n789), .B2(new_n273), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT99), .ZN(new_n863));
  INV_X1    g0663(.A(new_n781), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n861), .B(new_n863), .C1(G58), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n844), .B1(new_n845), .B2(new_n866), .C1(new_n830), .C2(new_n764), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n840), .A2(new_n867), .ZN(G384));
  NAND2_X1  g0668(.A1(new_n442), .A2(new_n440), .ZN(new_n869));
  INV_X1    g0669(.A(new_n441), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(G116), .A3(new_n217), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OR3_X1    g0675(.A1(new_n219), .A2(new_n267), .A3(new_n392), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n202), .A2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n253), .B(G13), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n405), .A2(new_n674), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n416), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n409), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n406), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n664), .A2(new_n881), .A3(new_n409), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n881), .B1(new_n413), .B2(new_n415), .ZN(new_n892));
  INV_X1    g0692(.A(new_n889), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT91), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n736), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(new_n724), .A3(new_n732), .A4(new_n731), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n719), .A2(new_n735), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n901), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT31), .B1(new_n901), .B2(new_n683), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(KEYINPUT106), .A3(new_n719), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n278), .A2(new_n675), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n662), .A2(new_n656), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n330), .B2(new_n335), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n831), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n880), .B1(new_n898), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n881), .B1(new_n665), .B2(new_n652), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n406), .A2(new_n885), .A3(new_n881), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n887), .A2(new_n922), .A3(KEYINPUT37), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n887), .A2(new_n922), .A3(KEYINPUT37), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n887), .B2(KEYINPUT37), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n886), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(KEYINPUT105), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n891), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n890), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(KEYINPUT40), .A3(new_n910), .A4(new_n915), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n917), .A2(G330), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n438), .A2(G330), .A3(new_n910), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT107), .Z(new_n937));
  AND2_X1   g0737(.A1(new_n917), .A2(new_n933), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n438), .A2(new_n910), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT39), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n662), .A2(new_n683), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n665), .A2(new_n674), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n896), .A2(new_n897), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n913), .A2(new_n914), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n434), .A2(new_n675), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n833), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n947), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n718), .A2(new_n438), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n668), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n940), .A2(new_n957), .B1(new_n253), .B2(new_n747), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n879), .B1(new_n959), .B2(new_n960), .ZN(G367));
  NOR2_X1   g0761(.A1(new_n522), .A2(new_n675), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n641), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n643), .A2(new_n683), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n685), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT42), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n965), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n572), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n675), .B1(new_n970), .B2(new_n712), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n683), .A2(new_n629), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n628), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n635), .B2(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n972), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n968), .A2(new_n971), .A3(new_n976), .A4(new_n975), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n700), .A2(new_n969), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n704), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n700), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n969), .B1(new_n688), .B2(new_n693), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n688), .A2(new_n693), .A3(new_n969), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n985), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n689), .ZN(new_n992));
  INV_X1    g0792(.A(G330), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n682), .B(new_n684), .C1(new_n698), .C2(new_n993), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n700), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n700), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n742), .B2(new_n744), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n986), .B(KEYINPUT45), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n989), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n700), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n991), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n984), .B1(new_n1003), .B2(new_n745), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n750), .A2(new_n253), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n983), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n766), .B1(new_n207), .B2(new_n428), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n236), .A2(new_n207), .A3(new_n371), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n752), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n789), .A2(new_n267), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n787), .A2(new_n340), .B1(new_n782), .B2(new_n223), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G68), .C2(new_n864), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n285), .B1(new_n774), .B2(new_n857), .C1(new_n777), .C2(new_n856), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n809), .B2(G50), .ZN(new_n1015));
  INV_X1    g0815(.A(G143), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1015), .C1(new_n798), .C2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n798), .A2(new_n851), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n371), .B1(new_n774), .B2(new_n1019), .C1(new_n777), .C2(new_n554), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n809), .B2(G283), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n804), .A2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n781), .A2(new_n419), .B1(new_n789), .B2(new_n225), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G303), .B2(new_n786), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1017), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1010), .B1(new_n1028), .B2(new_n762), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n975), .A2(new_n765), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1007), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT108), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT108), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1007), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1035), .ZN(G387));
  NOR2_X1   g0836(.A1(new_n998), .A2(new_n704), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n997), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n745), .B2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n755), .A2(new_n702), .B1(G107), .B2(new_n207), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n241), .A2(new_n451), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n702), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n339), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n759), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n752), .B1(new_n1047), .B2(new_n767), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n811), .A2(G159), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n771), .A2(new_n273), .B1(new_n774), .B2(new_n340), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n371), .B(new_n1050), .C1(new_n426), .C2(new_n854), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n789), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n786), .A2(G50), .B1(new_n1052), .B2(G97), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n864), .A2(new_n501), .B1(new_n804), .B2(G77), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n285), .B1(new_n775), .B2(G326), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n781), .A2(new_n790), .B1(new_n782), .B2(new_n554), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n786), .B1(new_n854), .B2(G311), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n783), .B2(new_n808), .C1(new_n798), .C2(new_n788), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1056), .B1(new_n583), .B2(new_n789), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1055), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1048), .B1(new_n1066), .B2(new_n762), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n682), .A2(new_n684), .A3(new_n765), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1038), .A2(new_n1006), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1039), .A2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n998), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n988), .A2(new_n990), .A3(new_n985), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n700), .B1(new_n999), .B2(new_n1001), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n751), .A3(new_n1003), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n797), .A2(new_n1019), .B1(new_n851), .B2(new_n787), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n285), .B1(new_n854), .B2(G303), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G294), .A2(new_n772), .B1(new_n775), .B2(G322), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n782), .A2(new_n790), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n813), .B(new_n1080), .C1(G116), .C2(new_n864), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n797), .A2(new_n340), .B1(new_n856), .B2(new_n787), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n781), .A2(new_n267), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n847), .B(new_n1085), .C1(G68), .C2(new_n804), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n285), .B1(new_n774), .B2(new_n1016), .C1(new_n777), .C2(new_n202), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n809), .B2(new_n426), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n845), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n766), .B1(new_n225), .B2(new_n207), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n249), .A2(new_n207), .A3(new_n371), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n752), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1090), .B(new_n1093), .C1(new_n969), .C2(new_n765), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n1006), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1075), .A2(new_n1096), .ZN(G390));
  AOI21_X1  g0897(.A(KEYINPUT106), .B1(new_n908), .B2(new_n719), .ZN(new_n1098));
  AND4_X1   g0898(.A1(KEYINPUT106), .A2(new_n719), .A3(new_n735), .A4(new_n902), .ZN(new_n1099));
  OAI211_X1 g0899(.A(G330), .B(new_n915), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT110), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT110), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n910), .A2(new_n1102), .A3(G330), .A4(new_n915), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n918), .B1(new_n929), .B2(KEYINPUT105), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n924), .A2(new_n925), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT38), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n890), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n943), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n945), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n833), .A2(new_n951), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n949), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1109), .A2(new_n941), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT109), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n912), .B1(new_n662), .B2(new_n656), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n330), .A2(new_n335), .A3(new_n911), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT109), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n675), .B(new_n830), .C1(new_n642), .C2(new_n715), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1118), .A2(new_n1119), .B1(new_n1120), .B2(new_n951), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1114), .A2(new_n1121), .A3(new_n945), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1104), .B1(new_n1113), .B2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1120), .A2(new_n951), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n932), .B(new_n1110), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n741), .A2(new_n830), .A3(new_n949), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n952), .A2(new_n945), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1127), .C1(new_n944), .C2(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1006), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n835), .B1(new_n841), .B2(new_n339), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n797), .A2(new_n1133), .B1(new_n860), .B2(new_n787), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT115), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n285), .B1(new_n789), .B2(new_n202), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT113), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n809), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n864), .A2(G159), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n854), .A2(G137), .B1(new_n775), .B2(G125), .ZN(new_n1143));
  AND4_X1   g0943(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n782), .A2(new_n340), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT53), .Z(new_n1147));
  NAND4_X1  g0947(.A1(new_n1135), .A2(new_n1137), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n811), .A2(G283), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n273), .A2(new_n789), .B1(new_n782), .B2(new_n373), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1085), .B(new_n1150), .C1(G116), .C2(new_n786), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n809), .A2(G97), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n371), .B1(new_n774), .B2(new_n554), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G107), .B2(new_n854), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1132), .B1(new_n845), .B2(new_n1156), .C1(new_n944), .C2(new_n764), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n950), .B1(new_n740), .B2(new_n831), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1101), .A2(new_n1103), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1111), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1127), .A2(new_n1125), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n910), .A2(G330), .A3(new_n830), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1124), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n935), .A2(new_n955), .A3(new_n668), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1165), .A2(new_n1129), .A3(new_n1123), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT111), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT111), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1166), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1130), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT112), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1130), .B2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(KEYINPUT112), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n751), .A3(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1131), .B(new_n1157), .C1(new_n1173), .C2(new_n1179), .ZN(G378));
  NAND2_X1  g0980(.A1(new_n343), .A2(new_n674), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n364), .B(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(new_n764), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n752), .B1(new_n842), .B2(G50), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n703), .B2(new_n371), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n789), .A2(new_n223), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n781), .A2(new_n273), .B1(new_n782), .B2(new_n267), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G107), .C2(new_n786), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n777), .A2(new_n225), .B1(new_n771), .B2(new_n428), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n703), .B(new_n371), .C1(new_n774), .C2(new_n790), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(new_n1194), .C1(new_n583), .C2(new_n797), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1188), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT118), .B(G124), .Z(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n775), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1140), .A2(new_n804), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n854), .A2(G132), .B1(new_n772), .B2(G137), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1133), .C2(new_n787), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n811), .A2(G125), .B1(G150), .B2(new_n864), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT117), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT117), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1199), .B1(new_n856), .B2(new_n789), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1197), .B1(new_n1196), .B2(new_n1195), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1186), .B1(new_n1211), .B2(new_n762), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1185), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1184), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n934), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n917), .A2(new_n1184), .A3(G330), .A4(new_n933), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1215), .A2(new_n954), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n954), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1213), .B1(new_n1219), .B2(new_n1005), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1167), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1219), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1168), .A2(KEYINPUT111), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1130), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1166), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n751), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1221), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT119), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(G375));
  OAI22_X1  g1032(.A1(new_n787), .A2(new_n790), .B1(new_n782), .B2(new_n225), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1011), .B(new_n1233), .C1(new_n501), .C2(new_n864), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n371), .B1(new_n774), .B2(new_n783), .C1(new_n777), .C2(new_n583), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n809), .B2(G107), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(new_n554), .C2(new_n797), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n787), .A2(new_n857), .B1(new_n782), .B2(new_n856), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1189), .B(new_n1238), .C1(G50), .C2(new_n864), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n811), .A2(G132), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1140), .A2(new_n854), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n285), .B1(new_n774), .B2(new_n1133), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G150), .B2(new_n772), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n845), .B1(new_n1237), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n835), .B(new_n1245), .C1(new_n273), .C2(new_n841), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT120), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1124), .B2(new_n763), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1165), .B2(new_n1006), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1171), .A2(new_n984), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1159), .A2(new_n1111), .B1(new_n1163), .B2(new_n1161), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1166), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1249), .B1(new_n1250), .B2(new_n1253), .ZN(G381));
  NAND2_X1  g1054(.A1(new_n1131), .A2(new_n1157), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1175), .A2(new_n751), .A3(new_n1178), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1039), .A2(new_n821), .A3(new_n1069), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G387), .A2(G381), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1231), .A2(new_n1258), .A3(new_n1264), .ZN(G407));
  NAND2_X1  g1065(.A1(new_n1231), .A2(new_n1258), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(new_n1266), .C2(G343), .ZN(G409));
  OAI211_X1 g1067(.A(G378), .B(new_n1221), .C1(new_n1224), .C2(new_n1229), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1227), .A2(new_n984), .A3(new_n1219), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1258), .B1(new_n1269), .B2(new_n1220), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G343), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G213), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT122), .B1(new_n840), .B2(new_n867), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT121), .B1(new_n1252), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT121), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1251), .A2(new_n1277), .A3(KEYINPUT60), .A4(new_n1166), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1252), .A2(new_n1275), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1171), .A2(new_n704), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1274), .B1(new_n1281), .B2(new_n1249), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n840), .A2(KEYINPUT122), .A3(new_n867), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(KEYINPUT122), .A3(new_n1260), .A4(new_n1249), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1271), .A2(new_n1273), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1283), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1274), .B(new_n1291), .C1(new_n1281), .C2(new_n1249), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1285), .ZN(new_n1293));
  INV_X1    g1093(.A(G2897), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n1292), .A2(new_n1293), .B1(new_n1294), .B2(new_n1273), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1273), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1284), .A2(G2897), .A3(new_n1296), .A4(new_n1285), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1286), .A3(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1289), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1007), .A2(G390), .A3(new_n1031), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT124), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n821), .B1(new_n1039), .B2(new_n1069), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1262), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT124), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1007), .A2(G390), .A3(new_n1309), .A4(new_n1031), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1305), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1033), .A2(new_n1035), .A3(new_n1259), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(KEYINPUT123), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1032), .A2(new_n1259), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT123), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1007), .A2(G390), .A3(new_n1315), .A4(new_n1031), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1311), .A2(new_n1312), .B1(new_n1317), .B2(new_n1307), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1303), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1271), .A2(new_n1273), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1317), .A2(new_n1307), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1328), .B1(new_n1300), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1287), .A2(new_n1321), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1320), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1318), .B1(new_n1300), .B2(new_n1322), .ZN(new_n1334));
  AND4_X1   g1134(.A1(new_n1320), .A2(new_n1299), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1319), .B1(new_n1333), .B2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(new_n1230), .A2(G378), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1266), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1318), .B(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1338), .B(new_n1340), .ZN(G402));
endmodule


