//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n462), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT69), .Z(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  MUX2_X1   g054(.A(G100), .B(G112), .S(G2105), .Z(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G2104), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n469), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT71), .Z(G162));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n462), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n468), .A2(new_n494), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT73), .A2(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT73), .A2(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n462), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n462), .A2(G102), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n479), .A2(KEYINPUT72), .A3(G126), .ZN(new_n502));
  OAI211_X1 g077(.A(G126), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n496), .A2(new_n501), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(G88), .A2(new_n511), .B1(new_n513), .B2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT5), .B(G543), .Z(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n526), .B(KEYINPUT77), .C1(new_n510), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n526), .B1(new_n510), .B2(new_n527), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(G63), .A3(G651), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(G90), .A2(new_n511), .B1(new_n513), .B2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n536), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n545), .A2(KEYINPUT78), .A3(G651), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT78), .B1(new_n545), .B2(G651), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n541), .B1(new_n546), .B2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n543), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n510), .A2(new_n554), .B1(new_n512), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  AOI22_X1  g142(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G651), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(G91), .B2(new_n511), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n508), .A2(KEYINPUT80), .A3(G53), .A4(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G166), .ZN(G303));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n569), .B1(new_n543), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n510), .A2(new_n578), .B1(new_n512), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n511), .A2(KEYINPUT83), .A3(G86), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n510), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n513), .A2(G48), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n509), .A2(new_n589), .A3(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n589), .B1(new_n509), .B2(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g171(.A(KEYINPUT82), .B(G651), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n588), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n543), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n569), .B1(new_n601), .B2(KEYINPUT84), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(KEYINPUT84), .B2(new_n601), .ZN(new_n603));
  AOI22_X1  g178(.A1(G85), .A2(new_n511), .B1(new_n513), .B2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n607));
  OR3_X1    g182(.A1(new_n510), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n510), .B2(new_n606), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n608), .B(new_n609), .C1(new_n569), .C2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n513), .A2(KEYINPUT86), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n512), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n612), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n618), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g194(.A(new_n618), .B(G301), .S(G868), .Z(G321));
  NOR2_X1   g195(.A1(G299), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g197(.A(new_n621), .B1(G168), .B2(G868), .ZN(G280));
  XNOR2_X1  g198(.A(KEYINPUT87), .B(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(G860), .B2(new_n624), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n560), .B(new_n626), .S(G868), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT88), .Z(G323));
  XOR2_X1   g203(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  INV_X1    g205(.A(new_n486), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G135), .ZN(new_n632));
  MUX2_X1   g207(.A(G99), .B(G111), .S(G2105), .Z(new_n633));
  AOI22_X1  g208(.A1(G123), .A2(new_n479), .B1(new_n633), .B2(G2104), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n484), .A2(G2104), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(KEYINPUT90), .B(KEYINPUT13), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n641), .A3(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  INV_X1    g220(.A(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2427), .ZN(new_n648));
  INV_X1    g223(.A(G2430), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT91), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n665), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT94), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n687), .B(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(G229));
  AND2_X1   g274(.A1(new_n462), .A2(G2104), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G103), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT98), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT25), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT99), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n462), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n631), .A2(G139), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n703), .B(new_n707), .C1(new_n704), .C2(new_n706), .ZN(new_n708));
  MUX2_X1   g283(.A(G33), .B(new_n708), .S(G29), .Z(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G2072), .Z(new_n710));
  NOR2_X1   g285(.A1(G4), .A2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n617), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1348), .Z(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NOR2_X1   g290(.A1(G168), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n715), .B2(G21), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n710), .B(new_n713), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n718), .B1(G2090), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G19), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n561), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT96), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G1341), .Z(new_n727));
  NOR2_X1   g302(.A1(new_n722), .A2(G2090), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n475), .B2(G29), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT100), .Z(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n719), .A2(G26), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  MUX2_X1   g315(.A(G104), .B(G116), .S(G2105), .Z(new_n741));
  AOI22_X1  g316(.A1(G128), .A2(new_n479), .B1(new_n741), .B2(G2104), .ZN(new_n742));
  INV_X1    g317(.A(G140), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n486), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT97), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2067), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n737), .A2(new_n738), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G105), .B2(new_n700), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n479), .A2(G129), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(new_n752), .C2(new_n751), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G141), .B2(new_n631), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G32), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(KEYINPUT102), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT102), .B2(new_n758), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT103), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n761), .A2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(G164), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G27), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n715), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n765), .A2(new_n766), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n715), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n715), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n717), .A2(new_n714), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT30), .A2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT30), .A2(G28), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT31), .B(G11), .Z(new_n783));
  INV_X1    g358(.A(new_n635), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(G29), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n779), .B(new_n785), .C1(new_n769), .C2(new_n768), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n775), .A2(new_n778), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n723), .A2(new_n729), .A3(new_n750), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n715), .A2(G23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n581), .B2(new_n715), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT33), .B(G1976), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(G303), .A2(G16), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n715), .A2(G22), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(G1971), .B1(new_n793), .B2(new_n794), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G6), .B(G305), .S(G16), .Z(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  XOR2_X1   g376(.A(new_n800), .B(new_n801), .Z(new_n802));
  OAI21_X1  g377(.A(KEYINPUT34), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT95), .Z(new_n804));
  NOR3_X1   g379(.A1(new_n799), .A2(KEYINPUT34), .A3(new_n802), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G24), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n603), .A2(new_n604), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G1986), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n631), .A2(G131), .ZN(new_n811));
  MUX2_X1   g386(.A(G95), .B(G107), .S(G2105), .Z(new_n812));
  AOI22_X1  g387(.A1(G119), .A2(new_n479), .B1(new_n812), .B2(G2104), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n805), .A2(new_n809), .A3(new_n810), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n804), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n788), .B1(new_n821), .B2(new_n823), .ZN(G311));
  INV_X1    g399(.A(new_n788), .ZN(new_n825));
  INV_X1    g400(.A(new_n823), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n822), .B1(new_n804), .B2(new_n819), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(G150));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G67), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n543), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G651), .ZN(new_n832));
  AOI22_X1  g407(.A1(G93), .A2(new_n511), .B1(new_n513), .B2(G55), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT104), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT105), .B(G860), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT107), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n617), .A2(G559), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT38), .Z(new_n844));
  NAND3_X1  g419(.A1(new_n835), .A2(new_n560), .A3(new_n837), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n561), .A2(new_n834), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n848), .A2(KEYINPUT106), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT106), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT108), .ZN(G145));
  XNOR2_X1  g430(.A(new_n475), .B(G162), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n784), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n631), .A2(G142), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT110), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(KEYINPUT111), .A3(G2105), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT111), .B1(new_n861), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n862), .A2(new_n865), .B1(new_n479), .B2(G130), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n814), .B(new_n638), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n493), .A2(new_n495), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n493), .B2(new_n495), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n745), .B(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n757), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n708), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n857), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(new_n878), .ZN(new_n886));
  INV_X1    g461(.A(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n857), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n885), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n882), .A2(new_n883), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT40), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n897), .ZN(G395));
  NOR2_X1   g473(.A1(new_n838), .A2(G868), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n847), .B(new_n626), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n617), .A2(G299), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT112), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n617), .A2(KEYINPUT112), .A3(G299), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n573), .B(new_n571), .C1(new_n611), .C2(new_n616), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n901), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(KEYINPUT41), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n905), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n902), .B2(new_n901), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n904), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(new_n900), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n807), .A2(new_n581), .ZN(new_n917));
  NAND2_X1  g492(.A1(G290), .A2(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G166), .A2(G305), .ZN(new_n920));
  OR2_X1    g495(.A1(G166), .A2(G305), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n917), .A3(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n915), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n915), .B2(new_n916), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n899), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n899), .B1(new_n928), .B2(G868), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(G301), .A2(G286), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(G301), .A2(G286), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n846), .B(new_n845), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n847), .A3(new_n933), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n938), .A3(new_n912), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT114), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n937), .A2(new_n847), .A3(new_n933), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n847), .B1(new_n933), .B2(new_n937), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT41), .B1(new_n911), .B2(new_n904), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n942), .A2(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT114), .A4(new_n912), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n932), .B1(new_n941), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n908), .B1(new_n942), .B2(new_n943), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n925), .A3(new_n939), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n953), .A2(new_n891), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n931), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n939), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n932), .ZN(new_n957));
  AND4_X1   g532(.A1(new_n931), .A2(new_n957), .A3(new_n891), .A4(new_n953), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT43), .B1(new_n951), .B2(new_n954), .ZN(new_n961));
  AND4_X1   g536(.A1(KEYINPUT43), .A2(new_n957), .A3(new_n891), .A4(new_n953), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n875), .B2(G1384), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n464), .A2(new_n465), .B1(new_n484), .B2(G137), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n471), .A2(new_n472), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(G40), .C1(new_n968), .C2(new_n462), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n745), .B(new_n748), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n757), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n972), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n975), .A2(KEYINPUT116), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(KEYINPUT116), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n970), .A2(new_n974), .B1(new_n978), .B2(new_n757), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n814), .A2(new_n817), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n748), .B2(new_n745), .ZN(new_n981));
  INV_X1    g556(.A(new_n970), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n816), .B1(new_n811), .B2(new_n813), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n970), .B1(new_n983), .B2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n970), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT48), .Z(new_n988));
  OAI22_X1  g563(.A1(new_n981), .A2(new_n982), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n978), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n976), .A2(KEYINPUT125), .A3(new_n990), .A4(new_n977), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n970), .B1(new_n971), .B2(new_n879), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n997));
  OR2_X1    g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n494), .B1(new_n484), .B2(G138), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT109), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n503), .B(KEYINPUT72), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(new_n501), .A3(new_n1004), .A4(new_n871), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n470), .A2(new_n473), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n581), .A2(G1976), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1010), .B1(G1976), .B2(new_n581), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n587), .B1(new_n510), .B2(new_n585), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1021), .B2(new_n594), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n588), .A2(new_n596), .A3(new_n1019), .A4(new_n597), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT120), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(KEYINPUT120), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT121), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1010), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1027), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1025), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1018), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n521), .A2(G8), .A3(new_n523), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n1038));
  XNOR2_X1  g613(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(KEYINPUT117), .B(KEYINPUT45), .C1(new_n506), .C2(new_n1008), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n493), .A2(new_n495), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1008), .B1(new_n873), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1044), .B2(new_n965), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n871), .A2(new_n501), .A3(new_n502), .A4(new_n505), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT45), .B(new_n1008), .C1(new_n1047), .C2(new_n874), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(new_n1007), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT50), .B(new_n1008), .C1(new_n1047), .C2(new_n874), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n969), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT118), .B(G2090), .Z(new_n1055));
  AOI22_X1  g630(.A1(new_n1050), .A2(new_n796), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1040), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1048), .A2(new_n1007), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1059), .A2(new_n1045), .A3(new_n1041), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G1971), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n969), .B1(new_n1044), .B2(KEYINPUT50), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1052), .B(new_n1008), .C1(new_n1047), .C2(new_n874), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1064), .A2(new_n1055), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1039), .B(G8), .C1(new_n1061), .C2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT45), .B(new_n1008), .C1(new_n873), .C2(new_n1043), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1067), .A2(new_n1007), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1966), .B1(new_n966), .B2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1062), .A2(new_n736), .A3(new_n1063), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G286), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1036), .A2(new_n1058), .A3(new_n1066), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1040), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1071), .A2(new_n1074), .A3(G286), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1036), .A2(new_n1077), .A3(new_n1066), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(new_n1013), .A3(new_n581), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1034), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1066), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1083), .A2(new_n1011), .B1(new_n1084), .B2(new_n1036), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1009), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1060), .B2(new_n972), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT59), .B1(new_n1090), .B2(new_n560), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1050), .B2(G1996), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n561), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT56), .B(G2072), .Z(new_n1097));
  NOR4_X1   g672(.A1(new_n1059), .A2(new_n1041), .A3(new_n1045), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1054), .A2(G1956), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G299), .B(KEYINPUT57), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n969), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1097), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1046), .A2(new_n1049), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1096), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1100), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT61), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1009), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n748), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(new_n618), .C1(new_n1064), .C2(G1348), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1348), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1009), .A2(G2067), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n617), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(KEYINPUT60), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1095), .A2(new_n1109), .A3(new_n1112), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1118), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1108), .B1(new_n1111), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1057), .B1(new_n533), .B2(new_n538), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1071), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT45), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1067), .A2(new_n1007), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n714), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1062), .A2(new_n736), .A3(new_n1063), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1057), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1137), .B2(new_n1127), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(G286), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1127), .B1(new_n1143), .B2(G8), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1144), .A2(new_n1131), .B1(G286), .B2(new_n1137), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(KEYINPUT123), .A3(new_n1138), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1050), .B2(G2078), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n966), .A2(new_n1068), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n769), .A2(KEYINPUT53), .ZN(new_n1151));
  OAI221_X1 g726(.A(new_n1149), .B1(G1961), .B2(new_n1064), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(G301), .B(KEYINPUT54), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n473), .A2(new_n1006), .A3(new_n1151), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(KEYINPUT124), .B2(new_n967), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(KEYINPUT124), .B2(new_n967), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1156), .A2(new_n966), .A3(new_n1048), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1064), .A2(G1961), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1153), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1152), .A2(new_n1153), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1126), .A2(new_n1147), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT123), .B1(new_n1145), .B2(new_n1138), .ZN(new_n1162));
  AND4_X1   g737(.A1(KEYINPUT123), .A2(new_n1132), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1142), .A2(new_n1146), .A3(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1152), .A2(G171), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1036), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1086), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(G290), .A2(KEYINPUT115), .A3(G1986), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT115), .ZN(new_n1173));
  INV_X1    g748(.A(G1986), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n807), .B2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n970), .B(new_n1172), .C1(new_n1175), .C2(new_n986), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n979), .A2(new_n984), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1000), .B1(new_n1171), .B2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g753(.A1(G227), .A2(new_n460), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1180), .A2(new_n661), .ZN(new_n1181));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n661), .A3(KEYINPUT127), .ZN(new_n1184));
  AOI21_X1  g758(.A(G229), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n885), .B2(new_n892), .ZN(new_n1186));
  NOR3_X1   g760(.A1(new_n1186), .A2(new_n961), .A3(new_n962), .ZN(G308));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n1188));
  OAI211_X1 g762(.A(new_n1188), .B(new_n1185), .C1(new_n885), .C2(new_n892), .ZN(G225));
endmodule


