//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NOR4_X1   g0018(.A1(new_n211), .A2(new_n214), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n203), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n225), .A2(new_n215), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n206), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n213), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n221), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n226), .A2(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n252), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n253), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(G238), .A3(new_n268), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n266), .A2(new_n275), .A3(new_n271), .A4(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT69), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n278), .A3(KEYINPUT13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G169), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(new_n282), .A3(G169), .A4(new_n279), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n274), .A2(G179), .A3(new_n276), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n230), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n267), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT12), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n292), .B2(new_n215), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n291), .A2(KEYINPUT12), .A3(G68), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n289), .A2(new_n215), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT65), .B1(G20), .B2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(KEYINPUT65), .A2(G20), .A3(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n231), .A2(G33), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n220), .B1(new_n222), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n231), .A2(G68), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n287), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n277), .A2(G200), .A3(new_n279), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n274), .A2(new_n276), .A3(G190), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n310), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT3), .B(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G238), .A2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(new_n226), .C2(G1698), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n265), .C1(G107), .C2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n264), .A2(new_n268), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G244), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n271), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G20), .A2(G77), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n324), .B1(new_n325), .B2(new_n300), .C1(new_n299), .C2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n287), .B1(new_n222), .B2(new_n292), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n222), .B2(new_n289), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n313), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  OAI21_X1  g0134(.A(G159), .B1(new_n297), .B2(new_n298), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G58), .A2(G68), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G58), .A2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(KEYINPUT70), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  INV_X1    g0141(.A(G159), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT65), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n231), .A3(new_n253), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(new_n296), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n231), .B1(new_n233), .B2(new_n336), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n255), .A2(KEYINPUT71), .A3(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n254), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n314), .B2(G20), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n215), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n334), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n257), .B2(new_n231), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n353), .B(G20), .C1(new_n254), .C2(new_n256), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n347), .A4(new_n340), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n287), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT64), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n326), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n225), .A2(KEYINPUT64), .A3(KEYINPUT8), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n289), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n292), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(G223), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n221), .A2(G1698), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n254), .A2(new_n371), .A3(new_n256), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(KEYINPUT73), .A3(new_n374), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n265), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n270), .B1(new_n319), .B2(G232), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(G190), .ZN(new_n382));
  AOI21_X1  g0182(.A(G200), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n363), .B(new_n369), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n384), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n373), .A2(KEYINPUT73), .A3(new_n374), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT73), .B1(new_n373), .B2(new_n374), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n390), .A2(new_n391), .A3(new_n264), .ZN(new_n392));
  INV_X1    g0192(.A(new_n380), .ZN(new_n393));
  OAI21_X1  g0193(.A(G169), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n381), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n363), .A2(KEYINPUT72), .A3(new_n369), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT72), .B1(new_n363), .B2(new_n369), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT18), .B(new_n396), .C1(new_n397), .C2(new_n398), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n389), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n258), .A2(G222), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n314), .B(new_n405), .C1(new_n370), .C2(new_n258), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n265), .C1(G77), .C2(new_n314), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n271), .C1(new_n221), .C2(new_n318), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G200), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n411));
  INV_X1    g0211(.A(G150), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n411), .B1(new_n412), .B2(new_n299), .C1(new_n367), .C2(new_n300), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n287), .B1(new_n220), .B2(new_n292), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n288), .A2(G50), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT9), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n409), .B1(new_n410), .B2(new_n408), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n416), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(KEYINPUT9), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT10), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT10), .B1(new_n418), .B2(new_n420), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n408), .A2(new_n330), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT66), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n408), .A2(G179), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n321), .ZN(new_n430));
  INV_X1    g0230(.A(G200), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n329), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT67), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(G190), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT67), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n432), .B2(new_n329), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n333), .A2(new_n404), .A3(new_n429), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT24), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n254), .A2(new_n256), .A3(new_n231), .A4(G87), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT22), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n314), .A2(KEYINPUT22), .A3(new_n231), .A4(G87), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT85), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n231), .B2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT23), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n447), .B(new_n450), .C1(new_n231), .C2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n445), .A2(new_n446), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n442), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n445), .A2(new_n446), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n453), .A4(new_n452), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(KEYINPUT24), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n287), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n267), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n291), .A2(new_n464), .A3(new_n230), .A4(new_n286), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT25), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n291), .B2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n469), .A2(G107), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n208), .A2(new_n258), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n210), .A2(G1698), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n314), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n265), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n267), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT77), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n267), .A4(G45), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n269), .B1(KEYINPUT5), .B2(new_n263), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n482), .A2(new_n486), .A3(new_n264), .A4(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n483), .A2(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n264), .B(G264), .C1(new_n481), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n480), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n431), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(G190), .B2(new_n491), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n463), .A2(new_n474), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  OAI21_X1  g0296(.A(G244), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n495), .A2(new_n497), .B1(KEYINPUT76), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n208), .A2(new_n258), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n314), .A2(new_n500), .B1(G33), .B2(G283), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n223), .B1(KEYINPUT76), .B2(new_n498), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n498), .A2(KEYINPUT76), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n314), .A2(new_n502), .A3(new_n258), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n265), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT78), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n264), .B(G257), .C1(new_n481), .C2(new_n489), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n488), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n506), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(G190), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n209), .A2(new_n472), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n472), .A2(KEYINPUT6), .A3(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G20), .ZN(new_n520));
  OAI21_X1  g0320(.A(G77), .B1(new_n297), .B2(new_n298), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n257), .A2(new_n231), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n520), .B(new_n521), .C1(new_n523), .C2(new_n472), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n287), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n291), .A2(G97), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n469), .B2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n506), .A2(new_n510), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n513), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n216), .A2(new_n258), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n223), .A2(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n254), .A2(new_n533), .A3(new_n256), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G116), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n264), .ZN(new_n540));
  INV_X1    g0340(.A(G45), .ZN(new_n541));
  OAI211_X1 g0341(.A(KEYINPUT79), .B(G250), .C1(new_n541), .C2(G1), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  AOI21_X1  g0343(.A(G274), .B1(new_n543), .B2(G250), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n267), .A2(G45), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n264), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT80), .B1(new_n546), .B2(new_n264), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(G200), .B1(new_n540), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n539), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n265), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n264), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n264), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n553), .A2(new_n558), .A3(G190), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n467), .A2(new_n468), .A3(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n325), .A2(new_n292), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n314), .A2(new_n231), .A3(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n516), .A2(new_n207), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n252), .A2(new_n231), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(KEYINPUT19), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n252), .B2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n287), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n560), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n550), .A2(new_n559), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n330), .B1(new_n540), .B2(new_n549), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n553), .A2(new_n558), .A3(new_n395), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n325), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n467), .A3(new_n468), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n561), .A3(new_n569), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n509), .B1(new_n265), .B2(new_n505), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n507), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n330), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n525), .A2(new_n527), .B1(new_n581), .B2(new_n395), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n494), .A2(new_n532), .A3(new_n579), .A4(new_n585), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n465), .A2(new_n212), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n292), .A2(new_n212), .ZN(new_n588));
  AOI21_X1  g0388(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n589));
  INV_X1    g0389(.A(G283), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n253), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n286), .A2(new_n230), .B1(G20), .B2(new_n212), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n591), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT20), .B1(new_n591), .B2(new_n592), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n587), .B(new_n588), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n264), .B1(new_n257), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G264), .A2(G1698), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n314), .B(new_n599), .C1(new_n210), .C2(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT83), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n264), .B(G270), .C1(new_n481), .C2(new_n489), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n488), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n488), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(G190), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n488), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT83), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n488), .A2(new_n602), .A3(new_n603), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n600), .B2(new_n598), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n596), .B(new_n606), .C1(new_n610), .C2(new_n431), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n595), .A2(G169), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(G179), .A3(new_n595), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(KEYINPUT21), .A3(G169), .A4(new_n595), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n611), .A2(new_n614), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  INV_X1    g0419(.A(new_n490), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n265), .B2(new_n479), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n330), .B1(new_n621), .B2(new_n488), .ZN(new_n622));
  AND4_X1   g0422(.A1(G179), .A2(new_n480), .A3(new_n488), .A4(new_n490), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n491), .A2(G169), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(G179), .A3(new_n488), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT86), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n463), .A2(new_n474), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n441), .A2(new_n586), .A3(new_n618), .A4(new_n628), .ZN(G372));
  MUX2_X1   g0429(.A(new_n385), .B(new_n388), .S(new_n384), .Z(new_n630));
  NOR2_X1   g0430(.A1(new_n332), .A2(new_n312), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n309), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n363), .A2(new_n369), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n396), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(new_n400), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n423), .B1(new_n427), .B2(new_n426), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n585), .A2(new_n494), .A3(new_n532), .A4(new_n579), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n463), .A2(new_n474), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n625), .A2(new_n626), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n578), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n583), .A2(new_n584), .A3(new_n578), .A4(new_n571), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n643), .B1(new_n641), .B2(new_n640), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT87), .B1(new_n586), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n646), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n637), .B1(new_n441), .B2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G20), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n267), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT88), .B(KEYINPUT27), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n640), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n624), .A2(new_n627), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n672), .A2(new_n674), .A3(new_n494), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n628), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n670), .A2(new_n596), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n643), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n618), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n642), .A2(new_n671), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n644), .A2(new_n671), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n204), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n516), .A2(new_n207), .A3(new_n212), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n267), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n695));
  INV_X1    g0495(.A(new_n691), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n694), .B(new_n695), .C1(new_n234), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT91), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n655), .A2(new_n670), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT95), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT95), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n655), .A2(new_n703), .A3(new_n670), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n651), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n648), .A2(new_n649), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n578), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n628), .A2(new_n643), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n586), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n670), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n532), .A2(new_n579), .A3(new_n585), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n628), .A2(new_n618), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(new_n494), .A4(new_n670), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n638), .A2(KEYINPUT94), .A3(new_n716), .A4(new_n670), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n553), .A2(new_n621), .A3(new_n558), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(G179), .A3(new_n610), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n511), .A2(new_n512), .B1(new_n722), .B2(KEYINPUT92), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(G179), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(KEYINPUT92), .B2(new_n722), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n580), .A2(new_n582), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n530), .A2(new_n491), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n553), .A2(new_n558), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n616), .A2(new_n734), .A3(new_n395), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n671), .B1(new_n732), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT31), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n742), .B(new_n671), .C1(new_n732), .C2(new_n739), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n719), .A2(new_n720), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n714), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n699), .B1(new_n747), .B2(G1), .ZN(G364));
  INV_X1    g0548(.A(new_n683), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n267), .B1(new_n659), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n691), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n682), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n230), .B1(G20), .B2(new_n330), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT99), .B(G317), .Z(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT33), .Z(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(new_n410), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n758), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n231), .B1(new_n766), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(G294), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n231), .A2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n431), .A2(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n231), .A2(new_n410), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n771), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n257), .B1(new_n772), .B2(new_n590), .C1(new_n597), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n770), .A2(new_n766), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G329), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n395), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n770), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n773), .A2(new_n781), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n779), .B1(new_n780), .B2(new_n782), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n774), .A2(new_n207), .ZN(new_n790));
  INV_X1    g0590(.A(new_n782), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G77), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n220), .B2(new_n763), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT32), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n776), .B2(new_n342), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n777), .A2(KEYINPUT32), .A3(G159), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n768), .A2(G97), .ZN(new_n798));
  INV_X1    g0598(.A(new_n772), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G107), .B1(G68), .B2(new_n760), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n257), .B1(new_n787), .B2(G58), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n756), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n752), .B(KEYINPUT96), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT97), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n755), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n247), .A2(G45), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n690), .A2(new_n314), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n541), .B2(new_n235), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n812), .A2(new_n815), .B1(new_n212), .B2(new_n690), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n314), .A2(G355), .A3(new_n204), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n803), .A2(new_n804), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n682), .B2(new_n808), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n754), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  AND4_X1   g0622(.A1(new_n329), .A2(new_n323), .A3(new_n331), .A4(new_n670), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n671), .A2(new_n329), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n438), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n332), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n701), .A2(new_n704), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n655), .A2(new_n670), .A3(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(new_n746), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n691), .B2(new_n751), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n257), .B1(new_n776), .B2(new_n780), .C1(new_n207), .C2(new_n772), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n798), .B1(new_n763), .B2(new_n597), .ZN(new_n834));
  INV_X1    g0634(.A(new_n774), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(G107), .C2(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n761), .A2(new_n590), .B1(new_n782), .B2(new_n212), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n838), .C1(new_n839), .C2(new_n788), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n782), .A2(new_n342), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n761), .A2(new_n412), .B1(new_n763), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n842), .B(new_n844), .C1(G143), .C2(new_n787), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n845), .A2(KEYINPUT34), .B1(new_n220), .B2(new_n774), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(KEYINPUT34), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n772), .A2(new_n215), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n768), .A2(G58), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n777), .A2(G132), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n847), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n852), .B2(new_n257), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n804), .B1(new_n853), .B2(new_n755), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n755), .A2(new_n805), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(G77), .B2(new_n856), .C1(new_n806), .C2(new_n826), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n832), .A2(new_n857), .ZN(G384));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n362), .A2(new_n287), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT70), .B1(new_n335), .B2(new_n339), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n345), .A2(new_n346), .A3(new_n341), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT16), .B1(new_n863), .B2(new_n361), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n369), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n396), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n669), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(new_n384), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n868), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT72), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n633), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n363), .A2(KEYINPUT72), .A3(new_n369), .ZN(new_n872));
  INV_X1    g0672(.A(new_n396), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n872), .B1(new_n873), .B2(new_n668), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n384), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT102), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n869), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n401), .A2(new_n402), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n867), .B1(new_n880), .B2(new_n630), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n859), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n669), .B1(new_n397), .B2(new_n398), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n399), .A2(new_n886), .A3(new_n875), .A4(new_n384), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n868), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(KEYINPUT38), .C1(new_n403), .C2(new_n867), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n384), .A3(new_n634), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n877), .B1(new_n892), .B2(KEYINPUT37), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n886), .B1(new_n630), .B2(new_n635), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n859), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT39), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n308), .A2(new_n671), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n635), .A2(new_n669), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n670), .A2(new_n306), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n901), .B(new_n312), .C1(new_n285), .C2(new_n307), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n308), .A2(new_n670), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n823), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n829), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n882), .A2(new_n890), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n900), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n705), .A2(new_n440), .A3(new_n713), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n637), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n909), .B(new_n911), .Z(new_n912));
  OAI21_X1  g0712(.A(new_n826), .B1(new_n902), .B2(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n719), .A2(new_n720), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n741), .A2(new_n743), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n890), .B2(new_n895), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n917), .A2(new_n918), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n744), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n440), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n890), .A2(new_n895), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT40), .B1(new_n907), .B2(new_n916), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(new_n745), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n440), .A2(new_n746), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n912), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n267), .B2(new_n659), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n212), .B1(new_n519), .B2(KEYINPUT35), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n232), .C1(KEYINPUT35), .C2(new_n519), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n336), .A2(G77), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n234), .A2(new_n934), .B1(G50), .B2(new_n215), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n658), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n930), .A2(new_n933), .A3(new_n936), .ZN(G367));
  OAI211_X1 g0737(.A(new_n532), .B(new_n585), .C1(new_n529), .C2(new_n670), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n671), .A2(new_n583), .A3(new_n584), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n688), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n688), .A2(new_n940), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n675), .A2(new_n687), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n678), .B2(new_n687), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT104), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n749), .B1(new_n948), .B2(KEYINPUT104), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n684), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n746), .B(new_n714), .C1(new_n946), .C2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n691), .B(new_n953), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n750), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n947), .A2(new_n938), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n585), .B1(new_n938), .B2(new_n674), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n670), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n670), .A2(new_n570), .ZN(new_n961));
  MUX2_X1   g0761(.A(new_n579), .B(new_n647), .S(new_n961), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n960), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n684), .A2(new_n940), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n955), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n804), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n243), .A2(new_n814), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n810), .B1(new_n204), .B2(new_n325), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT109), .B(G137), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n314), .B1(new_n776), .B2(new_n976), .C1(new_n788), .C2(new_n412), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n782), .A2(new_n220), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n767), .A2(new_n215), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n760), .A2(G159), .B1(new_n762), .B2(G143), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n225), .B2(new_n774), .C1(new_n222), .C2(new_n772), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n799), .A2(G97), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n774), .A2(new_n212), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n839), .B2(new_n761), .C1(KEYINPUT46), .C2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G303), .B2(new_n787), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT108), .B(G317), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n777), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT106), .B(G311), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n314), .B1(new_n762), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT107), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n988), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n782), .A2(new_n590), .B1(new_n767), .B2(new_n472), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT105), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n980), .A2(new_n982), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n972), .B1(new_n973), .B2(new_n974), .C1(new_n997), .C2(new_n756), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT110), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n808), .B2(new_n962), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n971), .A2(new_n1000), .ZN(G387));
  AOI22_X1  g0801(.A1(new_n787), .A2(G50), .B1(G150), .B2(new_n777), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n835), .A2(G77), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n575), .A2(new_n768), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n367), .A2(new_n761), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n983), .B1(new_n763), .B2(new_n342), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n314), .B1(new_n782), .B2(new_n215), .ZN(new_n1008));
  NOR4_X1   g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT112), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n787), .A2(new_n987), .B1(G303), .B2(new_n791), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n783), .B2(new_n763), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n760), .B2(new_n989), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT48), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n590), .B2(new_n767), .C1(new_n839), .C2(new_n774), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n257), .B1(new_n776), .B2(new_n764), .C1(new_n212), .C2(new_n772), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n804), .B1(new_n1019), .B2(new_n755), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n326), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n692), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(G68), .A2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT50), .B1(new_n326), .B2(G50), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1022), .A2(new_n541), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n813), .B(new_n1025), .C1(new_n240), .C2(new_n541), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n314), .A2(new_n692), .A3(new_n204), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G107), .C2(new_n204), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT111), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n811), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1020), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n679), .A2(new_n809), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1032), .A2(new_n1033), .B1(new_n751), .B2(new_n951), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n747), .A2(new_n951), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n691), .B1(new_n747), .B2(new_n951), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(G393));
  INV_X1    g0837(.A(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n946), .A2(new_n684), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n946), .A2(new_n684), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(KEYINPUT114), .A3(new_n1039), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1044), .A3(new_n751), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n787), .A2(G159), .B1(G150), .B2(new_n762), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n772), .A2(new_n207), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n314), .B1(new_n767), .B2(new_n222), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n774), .A2(new_n215), .B1(new_n782), .B2(new_n326), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n220), .B2(new_n761), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G143), .B2(new_n777), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT115), .Z(new_n1054));
  NOR2_X1   g0854(.A1(new_n782), .A2(new_n839), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n787), .A2(G311), .B1(G317), .B2(new_n762), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT116), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n761), .A2(new_n597), .B1(new_n772), .B2(new_n472), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n314), .B(new_n1059), .C1(G116), .C2(new_n768), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n783), .C2(new_n776), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1055), .B(new_n1061), .C1(G283), .C2(new_n835), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n755), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n810), .B1(new_n209), .B2(new_n204), .C1(new_n250), .C2(new_n814), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n938), .A2(new_n809), .A3(new_n939), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n972), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1045), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1035), .A2(new_n946), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n691), .C1(new_n1035), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(G390));
  AND2_X1   g0871(.A1(new_n787), .A2(G132), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n835), .A2(G150), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n768), .A2(G159), .ZN(new_n1075));
  INV_X1    g0875(.A(G125), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT54), .B(G143), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n776), .C1(new_n782), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(G128), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n314), .B1(new_n763), .B2(new_n1079), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1072), .A2(new_n1074), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n220), .B2(new_n772), .C1(new_n761), .C2(new_n976), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n763), .A2(new_n590), .B1(new_n767), .B2(new_n222), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n314), .B(new_n1083), .C1(new_n787), .C2(G116), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n791), .A2(G97), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n760), .A2(G107), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n848), .B(new_n790), .C1(G294), .C2(new_n777), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n756), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n804), .B(new_n1089), .C1(new_n367), .C2(new_n855), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n897), .B2(new_n806), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n825), .A2(new_n332), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n905), .B1(new_n711), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n904), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n898), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n923), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n891), .A2(new_n896), .B1(new_n906), .B2(new_n898), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1096), .A2(KEYINPUT117), .A3(new_n923), .A4(new_n1097), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n744), .A2(new_n745), .A3(new_n827), .A4(new_n904), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1104), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1091), .B1(new_n1108), .B2(new_n750), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n746), .A2(new_n826), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT118), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1095), .B1(new_n1111), .B2(new_n826), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1094), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n746), .B(new_n826), .C1(new_n1111), .C2(new_n1095), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n829), .A2(new_n905), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1095), .B1(new_n746), .B2(new_n826), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n1104), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n911), .A2(new_n927), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1105), .A2(new_n1107), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1122), .A2(new_n691), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1108), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1109), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G378));
  XOR2_X1   g0927(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n429), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n421), .A2(new_n422), .B1(new_n427), .B2(new_n426), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1128), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n419), .A2(new_n668), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1129), .A2(new_n1134), .A3(new_n1132), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT122), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(KEYINPUT122), .A3(new_n1137), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n805), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n763), .A2(new_n1076), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n788), .A2(new_n1079), .B1(new_n774), .B2(new_n1077), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G132), .C2(new_n760), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n843), .B2(new_n782), .C1(new_n412), .C2(new_n767), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT59), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(G33), .A2(G41), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT119), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G159), .B2(new_n799), .ZN(new_n1150));
  INV_X1    g0950(.A(G124), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n776), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n314), .A2(G41), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n220), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1147), .A2(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1003), .B1(new_n590), .B2(new_n776), .C1(new_n788), .C2(new_n472), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G58), .B2(new_n799), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n575), .A2(new_n791), .B1(G97), .B2(new_n760), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT120), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n979), .B1(new_n762), .B2(G116), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1153), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT58), .Z(new_n1162));
  OAI21_X1  g0962(.A(new_n755), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n752), .B1(new_n856), .B2(G50), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  NAND3_X1  g0965(.A1(new_n1142), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT123), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1137), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1134), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n926), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n926), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n917), .A2(new_n918), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n919), .A2(new_n916), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(KEYINPUT123), .A3(new_n1138), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1172), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n909), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n909), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1172), .A2(new_n1181), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1167), .B1(new_n1183), .B2(new_n751), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1180), .A2(new_n1182), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n691), .B1(new_n1185), .B2(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1122), .A2(new_n1121), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1184), .B1(new_n1186), .B2(new_n1188), .ZN(G375));
  OAI21_X1  g0989(.A(new_n314), .B1(new_n761), .B2(new_n1077), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n788), .A2(new_n976), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G132), .C2(new_n762), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n772), .A2(new_n225), .B1(new_n776), .B2(new_n1079), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G50), .B2(new_n768), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n412), .B2(new_n782), .C1(new_n342), .C2(new_n774), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1004), .B1(new_n788), .B2(new_n590), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT124), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n761), .A2(new_n212), .B1(new_n772), .B2(new_n222), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n314), .B(new_n1199), .C1(G294), .C2(new_n762), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n209), .B2(new_n774), .C1(new_n472), .C2(new_n782), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n776), .A2(new_n597), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n804), .B1(new_n1204), .B2(new_n755), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(G68), .B2(new_n856), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n904), .B2(new_n805), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1209));
  OAI211_X1 g1009(.A(KEYINPUT125), .B(new_n1208), .C1(new_n1209), .C2(new_n750), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n750), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1207), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n954), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT126), .ZN(G381));
  NAND2_X1  g1018(.A1(new_n1183), .A2(new_n751), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1166), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1168), .B(new_n1171), .C1(new_n920), .C2(G330), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT123), .B1(new_n1177), .B2(new_n1138), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1181), .B1(new_n1223), .B2(new_n1174), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1182), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1187), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n696), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1185), .A2(KEYINPUT57), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1220), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1126), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n971), .A2(new_n1067), .A3(new_n1070), .A4(new_n1000), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1231), .ZN(G409));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G375), .B2(G378), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n911), .A2(new_n927), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1209), .A2(new_n1241), .A3(KEYINPUT60), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1242), .A2(new_n1244), .A3(new_n691), .A4(new_n1124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n1214), .A3(G384), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1245), .B2(new_n1214), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1184), .B(new_n1126), .C1(new_n954), .C2(new_n1226), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n821), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1253), .A2(new_n1255), .A3(new_n1232), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1253), .B2(new_n1232), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1251), .A2(new_n1252), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT63), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1239), .A2(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1248), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1246), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT127), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1240), .A2(new_n1250), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(G2897), .A3(new_n1239), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1260), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G375), .A2(G378), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1239), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1249), .A3(new_n1271), .A4(new_n1250), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1259), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1271), .B(new_n1250), .C1(new_n1230), .C2(new_n1126), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1266), .A2(new_n1261), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1268), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1240), .A2(new_n1279), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(new_n1278), .A3(new_n1252), .A4(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1274), .A2(new_n1283), .ZN(G405));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1231), .A3(new_n1270), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1231), .A2(new_n1270), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1258), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1285), .A2(new_n1249), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1249), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


