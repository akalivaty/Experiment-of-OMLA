//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G113), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OR3_X1    g035(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT67), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n459), .B2(new_n460), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n466), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OR3_X1    g048(.A1(new_n466), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT68), .B1(new_n466), .B2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n466), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n483), .B2(G124), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n478), .A2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n482), .C1(new_n464), .C2(new_n465), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(G126), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n487), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n492));
  AND4_X1   g067(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(G164));
  NOR2_X1   g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT70), .B(G651), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT71), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n496), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n503), .A2(new_n504), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n507), .A2(G88), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n502), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND2_X1  g090(.A1(new_n507), .A2(G89), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT72), .B(G51), .Z(new_n517));
  NAND2_X1  g092(.A1(new_n500), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n521), .B1(new_n505), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n518), .A3(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G52), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n500), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n507), .A2(G90), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n496), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  NAND2_X1  g107(.A1(G68), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G56), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n510), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n508), .B1(new_n535), .B2(KEYINPUT74), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(KEYINPUT74), .B2(new_n535), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT75), .B(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n499), .B1(new_n506), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  INV_X1    g121(.A(G65), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n505), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n503), .A2(KEYINPUT79), .A3(new_n504), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT80), .B(G651), .C1(new_n551), .C2(new_n553), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(G91), .B2(new_n507), .ZN(new_n558));
  NAND2_X1  g133(.A1(G53), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT70), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT70), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT6), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n559), .B1(new_n564), .B2(new_n495), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT76), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n559), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n498), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n562), .A2(KEYINPUT70), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n560), .A2(G651), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n497), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n566), .B(new_n568), .C1(new_n575), .C2(new_n494), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n498), .A2(new_n578), .A3(new_n566), .A4(new_n568), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n572), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT78), .B1(new_n572), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n558), .B1(new_n581), .B2(new_n582), .ZN(G299));
  NAND2_X1  g158(.A1(new_n500), .A2(G49), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n507), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n505), .A2(G61), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(KEYINPUT81), .B1(G73), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n505), .A2(new_n590), .A3(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(new_n508), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n507), .A2(G86), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n500), .A2(G48), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n507), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n500), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n496), .C2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n507), .A2(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n549), .A2(new_n550), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n609), .A2(new_n562), .B1(new_n610), .B2(new_n499), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G284));
  XNOR2_X1  g188(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n556), .A2(new_n557), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n507), .A2(G91), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR3_X1   g194(.A1(new_n565), .A2(KEYINPUT76), .A3(new_n566), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n570), .B1(new_n569), .B2(KEYINPUT9), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n580), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n572), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n616), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n616), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n612), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n612), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n483), .A2(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n482), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n474), .A2(new_n475), .ZN(new_n638));
  INV_X1    g213(.A(G135), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n635), .B1(new_n636), .B2(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n482), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n640), .A2(G2096), .B1(new_n644), .B2(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n645), .B(new_n646), .C1(G2096), .C2(new_n640), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n654), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n655));
  AOI21_X1  g230(.A(KEYINPUT87), .B1(new_n654), .B2(KEYINPUT14), .ZN(new_n656));
  OAI22_X1  g231(.A1(new_n655), .A2(new_n656), .B1(new_n650), .B2(new_n653), .ZN(new_n657));
  XOR2_X1   g232(.A(G2443), .B(G2446), .Z(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(KEYINPUT88), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  INV_X1    g244(.A(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n676), .B1(new_n678), .B2(new_n674), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(new_n674), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT91), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n675), .A2(new_n676), .A3(new_n682), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n674), .A3(new_n676), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT18), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2096), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT92), .B(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XOR2_X1   g267(.A(G1971), .B(G1976), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n702), .B(new_n701), .S(new_n694), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n705), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n704), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(G229));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(G29), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n476), .A2(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G107), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n483), .B2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n717), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT94), .B(G16), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G24), .ZN(new_n731));
  INV_X1    g306(.A(G290), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n730), .ZN(new_n733));
  INV_X1    g308(.A(G1986), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n730), .A2(G22), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n730), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G6), .A2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G305), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT32), .B(G1981), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G23), .ZN(new_n746));
  INV_X1    g321(.A(G288), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n745), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT33), .B(G1976), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n739), .A2(new_n744), .A3(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n728), .B(new_n735), .C1(new_n751), .C2(KEYINPUT34), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(KEYINPUT34), .B2(new_n751), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT36), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n717), .A2(G35), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n717), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT29), .ZN(new_n757));
  INV_X1    g332(.A(G2090), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n730), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n541), .B2(new_n730), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT97), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1341), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G4), .A2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT95), .Z(new_n766));
  INV_X1    g341(.A(new_n612), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n745), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT96), .B(G1348), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n716), .A2(G26), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G128), .B2(new_n483), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n476), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n773), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT100), .B(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G11), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n782), .B1(new_n787), .B2(G28), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n786), .B1(new_n788), .B2(new_n789), .C1(new_n640), .C2(new_n716), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G34), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n716), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n472), .B2(new_n782), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n790), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n785), .B(new_n797), .C1(new_n791), .C2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n716), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n716), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G2078), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n782), .A2(G32), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n476), .A2(G141), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n470), .A2(G105), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT103), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n470), .A2(new_n806), .A3(G105), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n483), .A2(G129), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT26), .Z(new_n810));
  AND2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n802), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT27), .B(G1996), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n801), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n800), .A2(G2078), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n815), .B(new_n816), .C1(new_n813), .C2(new_n814), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n770), .A2(new_n798), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G127), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n466), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(G115), .A2(G2104), .ZN(new_n821));
  OAI21_X1  g396(.A(G2105), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT25), .Z(new_n824));
  INV_X1    g399(.A(G139), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n638), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT101), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT101), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  MUX2_X1   g404(.A(G33), .B(new_n829), .S(G29), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G2072), .ZN(new_n832));
  NAND2_X1  g407(.A1(G301), .A2(G16), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n745), .A2(G5), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G1961), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G168), .A2(new_n745), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n745), .B2(G21), .ZN(new_n839));
  INV_X1    g414(.A(G1966), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n839), .A2(new_n840), .B1(new_n836), .B2(new_n835), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n837), .B(new_n841), .C1(new_n840), .C2(new_n839), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n818), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n831), .A2(G2072), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n729), .A2(G20), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT23), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n626), .B2(new_n745), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1956), .ZN(new_n849));
  NOR4_X1   g424(.A1(new_n764), .A2(new_n843), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n754), .A2(new_n850), .ZN(G150));
  INV_X1    g426(.A(G150), .ZN(G311));
  OR2_X1    g427(.A1(new_n541), .A2(KEYINPUT106), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n541), .A2(KEYINPUT106), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n496), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT105), .ZN(new_n857));
  AOI22_X1  g432(.A1(G55), .A2(new_n500), .B1(new_n507), .B2(G93), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n859), .A2(new_n541), .A3(KEYINPUT106), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT38), .Z(new_n863));
  NOR2_X1   g438(.A1(new_n767), .A2(new_n629), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  NAND2_X1  g447(.A1(new_n483), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n482), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G142), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n638), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n642), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n725), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n829), .A2(KEYINPUT107), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n803), .A2(new_n811), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n803), .B2(new_n811), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n780), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n829), .A2(KEYINPUT107), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n781), .A3(new_n882), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n880), .A2(new_n885), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n829), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n879), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n891), .A3(new_n879), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n640), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(G162), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n889), .A2(new_n879), .A3(new_n891), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n892), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n902), .B2(new_n897), .ZN(new_n903));
  NOR4_X1   g478(.A1(new_n901), .A2(new_n892), .A3(new_n898), .A4(KEYINPUT108), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(G290), .B(G288), .ZN(new_n908));
  XNOR2_X1  g483(.A(G305), .B(KEYINPUT112), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G303), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n908), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(KEYINPUT113), .B2(KEYINPUT42), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT113), .B(KEYINPUT42), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n862), .B(new_n631), .Z(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n558), .B(new_n916), .C1(new_n581), .C2(new_n582), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n612), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n624), .A2(new_n625), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n919), .B2(new_n558), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n626), .A2(new_n916), .A3(new_n612), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G299), .A2(KEYINPUT110), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n612), .A3(new_n917), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n767), .A2(G299), .A3(KEYINPUT110), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT111), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n915), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n914), .A2(new_n924), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n914), .B1(new_n924), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n859), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n859), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  XOR2_X1   g516(.A(G286), .B(G301), .Z(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n862), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n929), .B2(new_n930), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n862), .B(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n923), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n911), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n933), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n934), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n911), .A3(new_n947), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n959));
  INV_X1    g534(.A(new_n923), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n944), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n931), .A2(new_n934), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n944), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n963), .B2(new_n911), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n946), .B1(new_n931), .B2(new_n934), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n949), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n941), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n965), .A3(new_n956), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n970), .A2(new_n959), .B1(new_n964), .B2(new_n950), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n941), .B2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n881), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n468), .A2(G40), .A3(new_n471), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n780), .A2(G2067), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n780), .A2(G2067), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n812), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n724), .B(new_n727), .Z(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n732), .A2(new_n734), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n732), .A2(new_n734), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n978), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n977), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n973), .A3(new_n881), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT116), .Z(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(G288), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n994), .B(new_n996), .C1(new_n995), .C2(G288), .ZN(new_n997));
  XNOR2_X1  g572(.A(G305), .B(G1981), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n994), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n993), .B(KEYINPUT116), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(G1976), .B2(new_n747), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n997), .B(new_n1000), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1007), .A2(KEYINPUT55), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(KEYINPUT55), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n977), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(KEYINPUT50), .B2(new_n974), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(G2090), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n976), .A2(new_n991), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n974), .A2(new_n975), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n738), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1012), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1013), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT117), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n1022));
  OR3_X1    g597(.A1(new_n974), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n758), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1012), .B1(new_n1025), .B2(new_n1018), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1005), .B(new_n1020), .C1(new_n1011), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1017), .ZN(new_n1028));
  INV_X1    g603(.A(G2078), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n991), .A4(new_n976), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT123), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1032), .A2(new_n1033), .B1(new_n836), .B2(new_n1014), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(KEYINPUT123), .A3(new_n1031), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1034), .A2(G301), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT125), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT124), .B(G2078), .Z(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1035), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1038), .A2(KEYINPUT125), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1049), .B(new_n1050), .C1(G171), .C2(new_n1043), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1040), .A2(G1966), .B1(new_n1014), .B2(G2084), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G168), .ZN(new_n1055));
  OAI21_X1  g630(.A(G8), .B1(new_n1053), .B2(G286), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(KEYINPUT51), .B2(new_n1056), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1040), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1024), .B2(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n558), .A2(new_n1063), .A3(new_n622), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1061), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1061), .A2(KEYINPUT121), .A3(new_n1065), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT61), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n992), .A2(G2067), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1014), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n612), .B1(new_n1076), .B2(KEYINPUT60), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT122), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1076), .A2(KEYINPUT60), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(new_n612), .C1(new_n1076), .C2(KEYINPUT60), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n541), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1040), .A2(new_n982), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n992), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT61), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1090), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1073), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1076), .A2(new_n767), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1067), .A2(new_n1068), .B1(new_n1097), .B2(new_n1092), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1052), .B(new_n1058), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1049), .B1(new_n1058), .B2(KEYINPUT62), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1054), .A2(new_n1012), .A3(G286), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1027), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1019), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1011), .B1(new_n1019), .B2(new_n1106), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1004), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1103), .B(new_n1020), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT63), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1000), .A2(new_n995), .A3(new_n747), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G1981), .B2(G305), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1020), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n994), .A2(new_n1115), .B1(new_n1005), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n990), .B1(new_n1105), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n978), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n986), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n987), .A2(new_n1120), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(KEYINPUT48), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(KEYINPUT48), .B2(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(new_n981), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n978), .B1(new_n1125), .B2(new_n812), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n978), .A2(new_n982), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT46), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT47), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n725), .A2(new_n727), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n979), .B1(new_n984), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n978), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1124), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g710(.A1(new_n970), .A2(new_n959), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n964), .A2(new_n950), .ZN(new_n1138));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g713(.A(G319), .ZN(new_n1140));
  NOR3_X1   g714(.A1(G229), .A2(G227), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n905), .A2(new_n672), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g716(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g717(.A(KEYINPUT126), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1145));
  AOI211_X1 g719(.A(new_n1145), .B(new_n1142), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1146));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1146), .ZN(G308));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n971), .B2(new_n1142), .ZN(new_n1148));
  NAND3_X1  g722(.A1(new_n1139), .A2(KEYINPUT126), .A3(new_n1143), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1149), .ZN(G225));
endmodule


