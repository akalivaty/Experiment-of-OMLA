

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U547 ( .A1(n677), .A2(G1384), .ZN(n767) );
  AND2_X2 U548 ( .A1(n515), .A2(G2104), .ZN(n862) );
  XNOR2_X1 U549 ( .A(n534), .B(KEYINPUT23), .ZN(n535) );
  BUF_X1 U550 ( .A(n691), .Z(n704) );
  INV_X1 U551 ( .A(n761), .ZN(n745) );
  INV_X1 U552 ( .A(n916), .ZN(n750) );
  INV_X1 U553 ( .A(G651), .ZN(n524) );
  BUF_X1 U554 ( .A(n540), .Z(n863) );
  NOR2_X2 U555 ( .A1(n622), .A2(n524), .ZN(n640) );
  NOR2_X2 U556 ( .A1(n544), .A2(n543), .ZN(G160) );
  XOR2_X1 U557 ( .A(n701), .B(KEYINPUT28), .Z(n510) );
  AND2_X1 U558 ( .A1(n919), .A2(n814), .ZN(n511) );
  AND2_X1 U559 ( .A1(n683), .A2(n682), .ZN(n684) );
  AND2_X1 U560 ( .A1(n685), .A2(n684), .ZN(n686) );
  INV_X1 U561 ( .A(n732), .ZN(n711) );
  NAND2_X1 U562 ( .A1(n711), .A2(G8), .ZN(n712) );
  OR2_X1 U563 ( .A1(n735), .A2(n712), .ZN(n713) );
  NOR2_X1 U564 ( .A1(n702), .A2(n510), .ZN(n703) );
  XNOR2_X1 U565 ( .A(n730), .B(n729), .ZN(n738) );
  NOR2_X2 U566 ( .A1(n767), .A2(n768), .ZN(n691) );
  INV_X1 U567 ( .A(n691), .ZN(n720) );
  NAND2_X1 U568 ( .A1(G8), .A2(n720), .ZN(n761) );
  NAND2_X1 U569 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U570 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n517) );
  NAND2_X1 U571 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U572 ( .A(KEYINPUT13), .ZN(n571) );
  NOR2_X1 U573 ( .A1(n801), .A2(n511), .ZN(n802) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n641) );
  XNOR2_X1 U575 ( .A(n536), .B(n535), .ZN(n538) );
  XNOR2_X1 U576 ( .A(n523), .B(n522), .ZN(n677) );
  BUF_X1 U577 ( .A(n677), .Z(G164) );
  AND2_X2 U578 ( .A1(G2104), .A2(G2105), .ZN(n866) );
  NAND2_X1 U579 ( .A1(G114), .A2(n866), .ZN(n513) );
  INV_X1 U580 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n515), .ZN(n539) );
  NAND2_X1 U582 ( .A1(G126), .A2(n539), .ZN(n512) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U584 ( .A(KEYINPUT88), .B(n514), .ZN(n521) );
  NAND2_X1 U585 ( .A1(G102), .A2(n862), .ZN(n519) );
  NOR2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n517), .B(n516), .ZN(n540) );
  NAND2_X1 U588 ( .A1(G138), .A2(n540), .ZN(n518) );
  NAND2_X1 U589 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U590 ( .A1(n521), .A2(n520), .ZN(n523) );
  INV_X1 U591 ( .A(KEYINPUT89), .ZN(n522) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n622) );
  NAND2_X1 U593 ( .A1(G78), .A2(n640), .ZN(n528) );
  NOR2_X1 U594 ( .A1(G543), .A2(n524), .ZN(n526) );
  XNOR2_X1 U595 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n525) );
  XNOR2_X2 U596 ( .A(n526), .B(n525), .ZN(n644) );
  NAND2_X1 U597 ( .A1(G65), .A2(n644), .ZN(n527) );
  NAND2_X1 U598 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U599 ( .A1(n641), .A2(G91), .ZN(n529) );
  XOR2_X1 U600 ( .A(KEYINPUT70), .B(n529), .Z(n530) );
  NOR2_X1 U601 ( .A1(n531), .A2(n530), .ZN(n533) );
  NOR2_X2 U602 ( .A1(G651), .A2(n622), .ZN(n645) );
  NAND2_X1 U603 ( .A1(n645), .A2(G53), .ZN(n532) );
  NAND2_X1 U604 ( .A1(n533), .A2(n532), .ZN(G299) );
  NAND2_X1 U605 ( .A1(G101), .A2(n862), .ZN(n536) );
  INV_X1 U606 ( .A(KEYINPUT64), .ZN(n534) );
  NAND2_X1 U607 ( .A1(G113), .A2(n866), .ZN(n537) );
  NAND2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n544) );
  BUF_X1 U609 ( .A(n539), .Z(n867) );
  NAND2_X1 U610 ( .A1(G125), .A2(n867), .ZN(n542) );
  NAND2_X1 U611 ( .A1(G137), .A2(n540), .ZN(n541) );
  NAND2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U613 ( .A1(G63), .A2(n644), .ZN(n546) );
  NAND2_X1 U614 ( .A1(G51), .A2(n645), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U616 ( .A(KEYINPUT6), .B(n547), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n641), .A2(G89), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U619 ( .A1(G76), .A2(n640), .ZN(n549) );
  NAND2_X1 U620 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U621 ( .A(n551), .B(KEYINPUT5), .Z(n552) );
  NOR2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U623 ( .A(KEYINPUT75), .B(n554), .Z(n555) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(n555), .Z(G168) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U626 ( .A(KEYINPUT9), .B(KEYINPUT69), .ZN(n559) );
  NAND2_X1 U627 ( .A1(G77), .A2(n640), .ZN(n557) );
  NAND2_X1 U628 ( .A1(G90), .A2(n641), .ZN(n556) );
  NAND2_X1 U629 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U630 ( .A(n559), .B(n558), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n645), .A2(G52), .ZN(n560) );
  XNOR2_X1 U632 ( .A(n560), .B(KEYINPUT68), .ZN(n562) );
  NAND2_X1 U633 ( .A1(G64), .A2(n644), .ZN(n561) );
  NAND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U635 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n565) );
  XOR2_X1 U640 ( .A(n565), .B(KEYINPUT10), .Z(n820) );
  NAND2_X1 U641 ( .A1(n820), .A2(G567), .ZN(n566) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  XOR2_X1 U643 ( .A(G860), .B(KEYINPUT72), .Z(n590) );
  NAND2_X1 U644 ( .A1(G56), .A2(n644), .ZN(n567) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n567), .Z(n574) );
  NAND2_X1 U646 ( .A1(n641), .A2(G81), .ZN(n568) );
  XNOR2_X1 U647 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U648 ( .A1(G68), .A2(n640), .ZN(n569) );
  NAND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U650 ( .A(n572), .B(n571), .ZN(n573) );
  NOR2_X1 U651 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n645), .A2(G43), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n924) );
  OR2_X1 U654 ( .A1(n590), .A2(n924), .ZN(G153) );
  XNOR2_X1 U655 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G79), .A2(n640), .ZN(n578) );
  NAND2_X1 U657 ( .A1(G54), .A2(n645), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U659 ( .A1(G66), .A2(n644), .ZN(n580) );
  NAND2_X1 U660 ( .A1(G92), .A2(n641), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U662 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U663 ( .A(n583), .B(KEYINPUT15), .Z(n606) );
  INV_X1 U664 ( .A(n606), .ZN(n922) );
  INV_X1 U665 ( .A(G868), .ZN(n659) );
  NAND2_X1 U666 ( .A1(n922), .A2(n659), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n584), .B(KEYINPUT74), .ZN(n586) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n586), .A2(n585), .ZN(G284) );
  XOR2_X1 U670 ( .A(KEYINPUT76), .B(G868), .Z(n587) );
  NOR2_X1 U671 ( .A1(G286), .A2(n587), .ZN(n589) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U673 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U674 ( .A1(G559), .A2(n590), .ZN(n591) );
  XOR2_X1 U675 ( .A(KEYINPUT77), .B(n591), .Z(n592) );
  NAND2_X1 U676 ( .A1(n592), .A2(n606), .ZN(n593) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n924), .ZN(n596) );
  NAND2_X1 U679 ( .A1(G868), .A2(n606), .ZN(n594) );
  NOR2_X1 U680 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U681 ( .A1(n596), .A2(n595), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n862), .ZN(n597) );
  XNOR2_X1 U683 ( .A(n597), .B(KEYINPUT78), .ZN(n600) );
  NAND2_X1 U684 ( .A1(G123), .A2(n867), .ZN(n598) );
  XNOR2_X1 U685 ( .A(n598), .B(KEYINPUT18), .ZN(n599) );
  NAND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U687 ( .A1(G111), .A2(n866), .ZN(n602) );
  NAND2_X1 U688 ( .A1(G135), .A2(n863), .ZN(n601) );
  NAND2_X1 U689 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n971) );
  XNOR2_X1 U691 ( .A(n971), .B(G2096), .ZN(n605) );
  INV_X1 U692 ( .A(G2100), .ZN(n825) );
  NAND2_X1 U693 ( .A1(n605), .A2(n825), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n606), .ZN(n607) );
  XNOR2_X1 U695 ( .A(n607), .B(n924), .ZN(n656) );
  NOR2_X1 U696 ( .A1(n656), .A2(G860), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G80), .A2(n640), .ZN(n609) );
  NAND2_X1 U698 ( .A1(G67), .A2(n644), .ZN(n608) );
  NAND2_X1 U699 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U700 ( .A1(G93), .A2(n641), .ZN(n610) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n610), .ZN(n611) );
  NOR2_X1 U702 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n645), .A2(G55), .ZN(n613) );
  NAND2_X1 U704 ( .A1(n614), .A2(n613), .ZN(n658) );
  XOR2_X1 U705 ( .A(n658), .B(KEYINPUT80), .Z(n615) );
  XNOR2_X1 U706 ( .A(n616), .B(n615), .ZN(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n645), .ZN(n618) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U709 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U710 ( .A(KEYINPUT81), .B(n619), .Z(n620) );
  NOR2_X1 U711 ( .A1(n644), .A2(n620), .ZN(n621) );
  XNOR2_X1 U712 ( .A(n621), .B(KEYINPUT82), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n622), .A2(G87), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U715 ( .A1(n645), .A2(G47), .ZN(n626) );
  NAND2_X1 U716 ( .A1(n644), .A2(G60), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U718 ( .A1(G72), .A2(n640), .ZN(n627) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n627), .Z(n628) );
  NOR2_X1 U720 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n641), .A2(G85), .ZN(n630) );
  NAND2_X1 U722 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U723 ( .A1(G73), .A2(n640), .ZN(n632) );
  XNOR2_X1 U724 ( .A(n632), .B(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U725 ( .A1(G61), .A2(n644), .ZN(n634) );
  NAND2_X1 U726 ( .A1(G86), .A2(n641), .ZN(n633) );
  NAND2_X1 U727 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U728 ( .A1(G48), .A2(n645), .ZN(n635) );
  XNOR2_X1 U729 ( .A(KEYINPUT83), .B(n635), .ZN(n636) );
  NOR2_X1 U730 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U731 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G75), .A2(n640), .ZN(n643) );
  NAND2_X1 U733 ( .A1(G88), .A2(n641), .ZN(n642) );
  NAND2_X1 U734 ( .A1(n643), .A2(n642), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G62), .A2(n644), .ZN(n647) );
  NAND2_X1 U736 ( .A1(G50), .A2(n645), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U738 ( .A1(n649), .A2(n648), .ZN(G166) );
  INV_X1 U739 ( .A(G166), .ZN(G303) );
  XOR2_X1 U740 ( .A(G290), .B(G305), .Z(n650) );
  XNOR2_X1 U741 ( .A(G288), .B(n650), .ZN(n651) );
  XOR2_X1 U742 ( .A(n651), .B(KEYINPUT19), .Z(n653) );
  XOR2_X1 U743 ( .A(G303), .B(KEYINPUT84), .Z(n652) );
  XNOR2_X1 U744 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U745 ( .A(n654), .B(G299), .ZN(n655) );
  XNOR2_X1 U746 ( .A(n655), .B(n658), .ZN(n891) );
  XNOR2_X1 U747 ( .A(n656), .B(n891), .ZN(n657) );
  NAND2_X1 U748 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U755 ( .A1(n665), .A2(G2072), .ZN(n666) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(n666), .Z(G158) );
  XNOR2_X1 U757 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G120), .A2(G69), .ZN(n667) );
  NOR2_X1 U760 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U761 ( .A1(G108), .A2(n668), .ZN(n912) );
  NAND2_X1 U762 ( .A1(n912), .A2(G567), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n669) );
  XNOR2_X1 U764 ( .A(KEYINPUT22), .B(n669), .ZN(n670) );
  NAND2_X1 U765 ( .A1(n670), .A2(G96), .ZN(n671) );
  NOR2_X1 U766 ( .A1(G218), .A2(n671), .ZN(n672) );
  XOR2_X1 U767 ( .A(KEYINPUT86), .B(n672), .Z(n913) );
  NAND2_X1 U768 ( .A1(n913), .A2(G2106), .ZN(n673) );
  NAND2_X1 U769 ( .A1(n674), .A2(n673), .ZN(n824) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n675) );
  XOR2_X1 U771 ( .A(KEYINPUT87), .B(n675), .Z(n676) );
  NOR2_X1 U772 ( .A1(n824), .A2(n676), .ZN(n823) );
  NAND2_X1 U773 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U774 ( .A1(G1348), .A2(n720), .ZN(n679) );
  NAND2_X1 U775 ( .A1(G2067), .A2(n704), .ZN(n678) );
  NAND2_X1 U776 ( .A1(n679), .A2(n678), .ZN(n688) );
  NOR2_X1 U777 ( .A1(n922), .A2(n688), .ZN(n687) );
  AND2_X1 U778 ( .A1(n704), .A2(G1996), .ZN(n681) );
  INV_X1 U779 ( .A(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U780 ( .A(n681), .B(n680), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n720), .A2(G1341), .ZN(n683) );
  INV_X1 U782 ( .A(n924), .ZN(n682) );
  NOR2_X1 U783 ( .A1(n687), .A2(n686), .ZN(n690) );
  AND2_X1 U784 ( .A1(n922), .A2(n688), .ZN(n689) );
  NOR2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n698) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n720), .ZN(n695) );
  INV_X1 U787 ( .A(KEYINPUT27), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n691), .A2(G2072), .ZN(n692) );
  XNOR2_X1 U789 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U791 ( .A(KEYINPUT95), .B(n696), .Z(n700) );
  NOR2_X1 U792 ( .A1(n700), .A2(G299), .ZN(n697) );
  NOR2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U794 ( .A(KEYINPUT96), .B(n699), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n700), .A2(G299), .ZN(n701) );
  XNOR2_X1 U796 ( .A(n703), .B(KEYINPUT29), .ZN(n708) );
  INV_X1 U797 ( .A(G1961), .ZN(n923) );
  NAND2_X1 U798 ( .A1(n720), .A2(n923), .ZN(n706) );
  XNOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .ZN(n993) );
  NAND2_X1 U800 ( .A1(n704), .A2(n993), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U802 ( .A1(G171), .A2(n709), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n719) );
  NOR2_X1 U804 ( .A1(G171), .A2(n709), .ZN(n710) );
  XOR2_X1 U805 ( .A(KEYINPUT97), .B(n710), .Z(n716) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n761), .ZN(n735) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n720), .ZN(n732) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n713), .ZN(n714) );
  NOR2_X1 U809 ( .A1(G168), .A2(n714), .ZN(n715) );
  NOR2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n717), .Z(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n731) );
  NAND2_X1 U813 ( .A1(n731), .A2(G286), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n761), .ZN(n722) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U817 ( .A(KEYINPUT99), .B(n723), .Z(n724) );
  NAND2_X1 U818 ( .A1(n724), .A2(G303), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT100), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n728), .A2(G8), .ZN(n730) );
  INV_X1 U822 ( .A(KEYINPUT32), .ZN(n729) );
  NAND2_X1 U823 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n731), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U826 ( .A(n736), .B(KEYINPUT98), .ZN(n737) );
  NOR2_X2 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U828 ( .A(n739), .B(KEYINPUT101), .ZN(n754) );
  NOR2_X1 U829 ( .A1(G288), .A2(G1976), .ZN(n740) );
  XOR2_X1 U830 ( .A(n740), .B(KEYINPUT102), .Z(n748) );
  INV_X1 U831 ( .A(n748), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n934) );
  NAND2_X1 U834 ( .A1(n754), .A2(n934), .ZN(n743) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n933) );
  NAND2_X1 U836 ( .A1(n743), .A2(n933), .ZN(n744) );
  XNOR2_X1 U837 ( .A(n744), .B(KEYINPUT103), .ZN(n746) );
  AND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n747), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n761), .A2(n748), .ZN(n749) );
  NAND2_X1 U841 ( .A1(KEYINPUT33), .A2(n749), .ZN(n751) );
  XNOR2_X1 U842 ( .A(G1981), .B(G305), .ZN(n916) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n765) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n754), .A2(n756), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n757), .B(KEYINPUT104), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n758), .A2(n761), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U850 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  OR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  INV_X1 U854 ( .A(n766), .ZN(n803) );
  INV_X1 U855 ( .A(n767), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n814) );
  XNOR2_X1 U857 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G104), .A2(n862), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G140), .A2(n863), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G116), .A2(n866), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G128), .A2(n867), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n779), .ZN(n888) );
  XNOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  NOR2_X1 U869 ( .A1(n888), .A2(n811), .ZN(n969) );
  NAND2_X1 U870 ( .A1(n814), .A2(n969), .ZN(n809) );
  INV_X1 U871 ( .A(n814), .ZN(n799) );
  NAND2_X1 U872 ( .A1(G107), .A2(n866), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G119), .A2(n867), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U875 ( .A(KEYINPUT91), .B(n782), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G95), .A2(n862), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G131), .A2(n863), .ZN(n783) );
  AND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n873) );
  NAND2_X1 U880 ( .A1(G1991), .A2(n873), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G105), .A2(n862), .ZN(n787) );
  XNOR2_X1 U882 ( .A(n787), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G129), .A2(n867), .ZN(n789) );
  NAND2_X1 U884 ( .A1(G141), .A2(n863), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n866), .A2(G117), .ZN(n790) );
  XOR2_X1 U887 ( .A(KEYINPUT92), .B(n790), .Z(n791) );
  NOR2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U890 ( .A(KEYINPUT93), .B(n795), .Z(n876) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n876), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT94), .B(n798), .Z(n984) );
  NOR2_X1 U894 ( .A1(n799), .A2(n984), .ZN(n806) );
  INV_X1 U895 ( .A(n806), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n809), .A2(n800), .ZN(n801) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n876), .ZN(n966) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n873), .ZN(n975) );
  NOR2_X1 U902 ( .A1(n804), .A2(n975), .ZN(n805) );
  NOR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n966), .A2(n807), .ZN(n808) );
  XNOR2_X1 U905 ( .A(KEYINPUT39), .B(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n888), .A2(n811), .ZN(n972) );
  NAND2_X1 U908 ( .A1(n812), .A2(n972), .ZN(n813) );
  XOR2_X1 U909 ( .A(KEYINPUT105), .B(n813), .Z(n815) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n819) );
  XNOR2_X1 U912 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n819), .B(n818), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n820), .ZN(G217) );
  INV_X1 U915 ( .A(n820), .ZN(G223) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U917 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U920 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U921 ( .A(n824), .ZN(G319) );
  XNOR2_X1 U922 ( .A(n825), .B(G2096), .ZN(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT42), .B(G2678), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT43), .B(G2090), .Z(n829) );
  XNOR2_X1 U926 ( .A(G2067), .B(G2072), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U929 ( .A(G2078), .B(G2084), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(G227) );
  XNOR2_X1 U931 ( .A(G1981), .B(n923), .ZN(n836) );
  INV_X1 U932 ( .A(G1996), .ZN(n834) );
  XOR2_X1 U933 ( .A(n834), .B(G1986), .Z(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U935 ( .A(G1976), .B(G1971), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1956), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U938 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2474), .B(KEYINPUT41), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1991), .B(KEYINPUT109), .Z(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U943 ( .A1(n867), .A2(G124), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U945 ( .A1(G100), .A2(n862), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U947 ( .A1(G112), .A2(n866), .ZN(n849) );
  NAND2_X1 U948 ( .A1(G136), .A2(n863), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U950 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G118), .A2(n866), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G130), .A2(n867), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n860) );
  NAND2_X1 U954 ( .A1(n862), .A2(G106), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT110), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G142), .A2(n863), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT45), .B(n857), .ZN(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(n858), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(G164), .B(n861), .ZN(n887) );
  XNOR2_X1 U962 ( .A(G162), .B(n971), .ZN(n875) );
  NAND2_X1 U963 ( .A1(G103), .A2(n862), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G139), .A2(n863), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n872) );
  NAND2_X1 U966 ( .A1(G115), .A2(n866), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G127), .A2(n867), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n978) );
  XNOR2_X1 U971 ( .A(n873), .B(n978), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT116), .B(KEYINPUT112), .ZN(n878) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT48), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(n880), .B(n879), .Z(n885) );
  XOR2_X1 U977 ( .A(KEYINPUT115), .B(KEYINPUT113), .Z(n882) );
  XNOR2_X1 U978 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(G160), .B(n883), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U984 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U985 ( .A(G286), .B(n891), .ZN(n893) );
  XOR2_X1 U986 ( .A(n924), .B(n922), .Z(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n895) );
  XNOR2_X1 U988 ( .A(G171), .B(KEYINPUT117), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2454), .B(G2435), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2438), .B(G2427), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n905) );
  XOR2_X1 U994 ( .A(KEYINPUT107), .B(G2446), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2443), .B(G2430), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n901), .B(G2451), .Z(n903) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(n906), .A2(G14), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n914), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  XOR2_X1 U1008 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1010 ( .A(G120), .ZN(G236) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(G325) );
  INV_X1 U1014 ( .A(G325), .ZN(G261) );
  INV_X1 U1015 ( .A(n914), .ZN(G401) );
  XOR2_X1 U1016 ( .A(KEYINPUT56), .B(G16), .Z(n939) );
  XOR2_X1 U1017 ( .A(G168), .B(G1966), .Z(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1019 ( .A(KEYINPUT57), .B(n917), .Z(n932) );
  XNOR2_X1 U1020 ( .A(G1956), .B(G299), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(G1971), .A2(G303), .ZN(n920) );
  NAND2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n930) );
  XOR2_X1 U1024 ( .A(n922), .B(G1348), .Z(n928) );
  XNOR2_X1 U1025 ( .A(G171), .B(n923), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n924), .B(G1341), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT125), .B(n937), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT126), .ZN(n964) );
  XOR2_X1 U1036 ( .A(G1966), .B(G21), .Z(n942) );
  XOR2_X1 U1037 ( .A(G1961), .B(G5), .Z(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n952) );
  XOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .Z(n943) );
  XNOR2_X1 U1040 ( .A(G4), .B(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G20), .B(G1956), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1341), .B(G19), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT60), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G1986), .B(KEYINPUT127), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(G24), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT58), .B(n958), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT61), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n962), .A2(G16), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n992) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT51), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n977) );
  XOR2_X1 U1064 ( .A(G2084), .B(G160), .Z(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n986) );
  XNOR2_X1 U1069 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G2072), .B(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G164), .B(G2078), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n982), .B(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT52), .B(n987), .Z(n988) );
  NOR2_X1 U1077 ( .A1(KEYINPUT55), .A2(n988), .ZN(n989) );
  XOR2_X1 U1078 ( .A(KEYINPUT120), .B(n989), .Z(n990) );
  NAND2_X1 U1079 ( .A1(G29), .A2(n990), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n1018) );
  XNOR2_X1 U1081 ( .A(n993), .B(G27), .ZN(n995) );
  XOR2_X1 U1082 ( .A(G1996), .B(G32), .Z(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n996), .ZN(n1002) );
  XOR2_X1 U1085 ( .A(G2067), .B(G26), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n997), .A2(G28), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(G2072), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G33), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G25), .B(G1991), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT53), .B(n1005), .Z(n1008) );
  XOR2_X1 U1094 ( .A(KEYINPUT54), .B(G34), .Z(n1006) );
  XNOR2_X1 U1095 ( .A(G2084), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(KEYINPUT121), .B(G2090), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(G35), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT55), .ZN(n1014) );
  INV_X1 U1101 ( .A(G29), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(G11), .A2(n1015), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT124), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1019), .Z(G150) );
  INV_X1 U1107 ( .A(G150), .ZN(G311) );
endmodule

