//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(G20), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n221), .B1(new_n202), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G58), .B2(G232), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT64), .B(G77), .Z(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G244), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n219), .A2(new_n220), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n209), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n215), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n206), .B2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT12), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n253), .B1(new_n255), .B2(new_n252), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n251), .A2(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n207), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n260), .B1(new_n207), .B2(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n263), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT11), .B1(new_n263), .B2(new_n249), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  OAI211_X1 g0073(.A(G226), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G97), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n285), .B2(G238), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT13), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT13), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n280), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n269), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n268), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  INV_X1    g0094(.A(new_n290), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n280), .B2(new_n286), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n293), .A2(KEYINPUT14), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n292), .B(G169), .C1(new_n295), .C2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n291), .A2(new_n268), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n267), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n267), .B1(new_n297), .B2(G190), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n297), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G222), .A2(G1698), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n273), .A2(G223), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n279), .C1(new_n225), .C2(new_n310), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n282), .B1(new_n285), .B2(G226), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n294), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n254), .A2(G50), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n250), .B2(G50), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT67), .ZN(new_n321));
  INV_X1    g0121(.A(G58), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(KEYINPUT8), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT8), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT67), .A3(G58), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(KEYINPUT8), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(G20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n249), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n320), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n316), .A2(new_n269), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n318), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n334), .B(KEYINPUT9), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n317), .A2(G190), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n307), .C2(new_n317), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n251), .A2(new_n261), .B1(new_n225), .B2(new_n254), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n324), .A2(G58), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n326), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n259), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  INV_X1    g0147(.A(new_n225), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n346), .B1(new_n262), .B2(new_n347), .C1(new_n348), .C2(new_n207), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n249), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n310), .A2(G232), .A3(new_n273), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n310), .A2(G238), .A3(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G107), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n310), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n279), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n282), .B1(new_n285), .B2(G244), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n357), .B2(new_n269), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n294), .A3(new_n356), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n350), .C1(new_n362), .C2(new_n357), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n309), .A2(new_n342), .A3(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(KEYINPUT3), .A2(G33), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT3), .A2(G33), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n270), .A2(new_n271), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n310), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G68), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n322), .A2(new_n252), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n201), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n259), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n252), .B1(new_n374), .B2(new_n368), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n380), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n385), .A3(new_n249), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n327), .A2(new_n254), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n250), .B2(new_n327), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(G223), .A2(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n222), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(new_n270), .C2(new_n271), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n278), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G232), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n281), .B1(new_n284), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT71), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n394), .B2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n269), .B1(new_n294), .B2(new_n397), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n389), .A2(KEYINPUT18), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT72), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n389), .A2(new_n402), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI211_X1 g0207(.A(KEYINPUT72), .B(KEYINPUT18), .C1(new_n389), .C2(new_n402), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n282), .B1(new_n285), .B2(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n392), .A2(new_n393), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n279), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT71), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n307), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n397), .A2(new_n362), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n386), .A3(new_n388), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n388), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n380), .B1(new_n375), .B2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n333), .B1(new_n422), .B2(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n385), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n417), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n409), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT80), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G294), .ZN(new_n429));
  INV_X1    g0229(.A(G294), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  OAI21_X1  g0231(.A(G33), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n433));
  OAI211_X1 g0233(.A(G250), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n279), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT5), .B(G41), .ZN(new_n437));
  INV_X1    g0237(.A(G45), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(G1), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n437), .A2(G274), .A3(new_n278), .A4(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n437), .A2(new_n439), .B1(new_n216), .B2(new_n277), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G264), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n307), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n435), .A2(new_n279), .B1(new_n441), .B2(G264), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n362), .A3(new_n440), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n207), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n310), .A2(new_n450), .A3(new_n207), .A4(G87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n207), .B2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n353), .A2(KEYINPUT23), .A3(G20), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n452), .A2(new_n453), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n452), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n249), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n254), .A2(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT79), .B(KEYINPUT25), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n206), .A2(G33), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n333), .A2(new_n254), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n353), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n443), .A2(new_n470), .A3(new_n307), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n447), .A2(new_n462), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n443), .A2(new_n269), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n445), .A2(new_n294), .A3(new_n440), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n452), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n452), .A2(new_n453), .A3(new_n459), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n333), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n469), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n473), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n374), .A2(new_n368), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G107), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n259), .A2(G77), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g0285(.A(G97), .B(G107), .Z(new_n486));
  INV_X1    g0286(.A(KEYINPUT6), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT73), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT6), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT74), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(new_n492), .C1(G97), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(G97), .B(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n495), .A3(new_n491), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n207), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n249), .B1(new_n485), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n254), .A2(G97), .ZN(new_n499));
  INV_X1    g0299(.A(new_n467), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G97), .ZN(new_n501));
  OAI211_X1 g0301(.A(G244), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G250), .A2(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(KEYINPUT4), .A2(G244), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G1698), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n310), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n278), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n439), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n278), .ZN(new_n515));
  INV_X1    g0315(.A(G257), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n440), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(G200), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n511), .A2(new_n517), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G190), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n498), .A2(new_n501), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n269), .B1(new_n511), .B2(new_n517), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n294), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n482), .A2(G107), .B1(G77), .B2(new_n259), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n486), .A2(new_n492), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n493), .A2(G97), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n496), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n333), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n501), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n522), .B(new_n523), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n521), .A2(new_n531), .A3(KEYINPUT75), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n481), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n500), .A2(G116), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n255), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n505), .B(new_n207), .C1(G33), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n249), .C1(new_n207), .C2(G116), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n537), .B(new_n539), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n206), .A2(G45), .ZN(new_n547));
  INV_X1    g0347(.A(new_n513), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT5), .A2(G41), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G274), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n216), .B2(new_n277), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n441), .A2(G270), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n366), .A2(G303), .A3(new_n367), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n279), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n546), .A2(new_n559), .A3(G169), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n553), .A2(G179), .A3(new_n558), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n560), .A2(new_n561), .B1(new_n546), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n553), .A2(new_n558), .A3(G190), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n546), .B1(G200), .B2(new_n559), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n310), .A2(KEYINPUT76), .A3(G238), .A4(new_n273), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n310), .A2(G244), .A3(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n454), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n279), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n547), .A2(G250), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n278), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n551), .B2(new_n547), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n269), .ZN(new_n581));
  XOR2_X1   g0381(.A(new_n347), .B(KEYINPUT77), .Z(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n500), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n310), .A2(new_n207), .A3(G68), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n207), .B1(new_n275), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n540), .A3(new_n353), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n585), .B1(new_n262), .B2(new_n540), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n249), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n347), .A2(new_n255), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n581), .B(new_n594), .C1(G179), .C2(new_n580), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n580), .A2(new_n362), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n500), .A2(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n598), .A3(new_n593), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n580), .B2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT78), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n578), .B1(new_n574), .B2(new_n279), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n307), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT78), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n536), .A2(new_n568), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n365), .A2(new_n427), .A3(new_n607), .ZN(G372));
  INV_X1    g0408(.A(new_n336), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n420), .A2(new_n425), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n308), .A2(new_n359), .A3(new_n358), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n305), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n613), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n269), .B1(new_n413), .B2(new_n414), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n397), .A2(new_n294), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n406), .B1(new_n424), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n403), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n340), .A2(new_n341), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n609), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n365), .A2(new_n427), .ZN(new_n624));
  INV_X1    g0424(.A(new_n531), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n600), .B1(new_n362), .B2(new_n580), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n595), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n595), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n602), .A2(new_n605), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n595), .A3(new_n625), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT82), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n480), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n462), .A2(new_n469), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(KEYINPUT82), .A3(new_n473), .A4(new_n474), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n565), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n626), .A2(new_n595), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n521), .A2(new_n531), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n472), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n630), .B(new_n633), .C1(new_n638), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n624), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(new_n643), .ZN(G369));
  INV_X1    g0444(.A(G330), .ZN(new_n645));
  INV_X1    g0445(.A(new_n546), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n568), .B1(new_n646), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n565), .A2(new_n546), .A3(new_n652), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n636), .A2(new_n652), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n472), .A2(new_n480), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT84), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT84), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n472), .A2(new_n657), .A3(new_n480), .A4(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n659), .B(new_n661), .C1(new_n480), .C2(new_n653), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n635), .A2(new_n637), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n652), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n565), .A2(new_n653), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n210), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n588), .A2(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n213), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n519), .A2(G179), .ZN(new_n679));
  AND4_X1   g0479(.A1(new_n580), .A2(new_n679), .A3(new_n559), .A4(new_n443), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT85), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n563), .A2(new_n603), .A3(new_n445), .A4(new_n519), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n603), .A2(new_n445), .A3(new_n519), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(KEYINPUT85), .A3(KEYINPUT30), .A4(new_n563), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n680), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n603), .A2(new_n519), .A3(new_n445), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n553), .A2(new_n558), .A3(G179), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n678), .B(new_n653), .C1(new_n687), .C2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n686), .ZN(new_n693));
  INV_X1    g0493(.A(new_n680), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n682), .A2(KEYINPUT86), .A3(new_n683), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT86), .B1(new_n682), .B2(new_n683), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n652), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT87), .B1(new_n700), .B2(new_n678), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT86), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n690), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n696), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n653), .B1(new_n687), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT87), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT31), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n692), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n700), .A2(KEYINPUT87), .A3(new_n678), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n706), .B1(new_n705), .B2(KEYINPUT31), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n691), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n536), .A2(new_n568), .A3(new_n606), .A4(new_n653), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT89), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n595), .A2(new_n640), .A3(new_n472), .A4(new_n626), .ZN(new_n718));
  INV_X1    g0518(.A(new_n565), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n664), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n629), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n652), .B1(new_n721), .B2(new_n633), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n717), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n625), .A2(new_n626), .A3(new_n595), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n596), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n631), .A2(new_n627), .A3(new_n595), .A4(new_n625), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n480), .A2(new_n562), .A3(new_n564), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n725), .B(new_n726), .C1(new_n641), .C2(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT29), .B1(new_n642), .B2(new_n653), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(KEYINPUT89), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n716), .A2(G330), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n677), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(new_n656), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n654), .A2(new_n645), .A3(new_n655), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n207), .A2(G13), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n206), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n672), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n654), .A2(new_n655), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n210), .A2(new_n310), .ZN(new_n746));
  INV_X1    g0546(.A(G355), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n210), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n671), .A2(new_n310), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n438), .B2(new_n214), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n243), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n215), .B1(G20), .B2(new_n269), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n744), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n739), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(new_n362), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n307), .A2(G179), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n587), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(G179), .A3(new_n307), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n294), .A2(new_n307), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n322), .B1(new_n765), .B2(new_n202), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n762), .B(new_n766), .C1(G107), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n767), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n310), .B1(new_n771), .B2(new_n252), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G97), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n767), .A2(new_n773), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n767), .A2(G179), .A3(new_n307), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n225), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n770), .A2(new_n776), .A3(new_n780), .A4(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n771), .A2(new_n788), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n765), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n310), .B(new_n790), .C1(G326), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n763), .ZN(new_n793));
  INV_X1    g0593(.A(new_n761), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(G322), .B1(new_n794), .B2(G303), .ZN(new_n795));
  INV_X1    g0595(.A(new_n777), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G283), .A2(new_n769), .B1(new_n796), .B2(G329), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n429), .A2(new_n431), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n775), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n792), .A2(new_n795), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n787), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n754), .B1(new_n803), .B2(KEYINPUT92), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n745), .B(new_n758), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n741), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  INV_X1    g0608(.A(new_n715), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n708), .B2(new_n709), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n645), .B1(new_n810), .B2(new_n714), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n363), .B1(new_n350), .B2(new_n653), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n360), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n358), .A2(new_n359), .A3(new_n653), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT93), .Z(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  MUX2_X1   g0617(.A(new_n816), .B(new_n817), .S(new_n722), .Z(new_n818));
  NOR2_X1   g0618(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT94), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT94), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n739), .B1(new_n811), .B2(new_n818), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n754), .A2(new_n742), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n740), .B1(new_n261), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n754), .ZN(new_n826));
  INV_X1    g0626(.A(new_n771), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G107), .A2(new_n794), .B1(new_n827), .B2(G283), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n789), .B2(new_n777), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n768), .A2(new_n587), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G294), .B2(new_n793), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n310), .B1(new_n791), .B2(G303), .ZN(new_n832));
  INV_X1    g0632(.A(new_n775), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n832), .C1(new_n540), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n829), .B(new_n834), .C1(G116), .C2(new_n785), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n793), .A2(G143), .B1(new_n791), .B2(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n771), .C1(new_n784), .C2(new_n778), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G50), .A2(new_n794), .B1(new_n796), .B2(G132), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n370), .B1(new_n769), .B2(G68), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n322), .C2(new_n833), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n835), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n825), .B1(new_n826), .B2(new_n845), .C1(new_n815), .C2(new_n743), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n823), .A2(new_n846), .ZN(G384));
  OR2_X1    g0647(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n215), .A2(new_n207), .A3(new_n538), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT95), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n348), .A2(new_n213), .A3(new_n377), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n202), .B2(G68), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n855), .A2(new_n206), .A3(G13), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT96), .ZN(new_n857));
  INV_X1    g0657(.A(new_n305), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n653), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n382), .A2(new_n249), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n422), .A2(KEYINPUT16), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n388), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n650), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n409), .B2(new_n426), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n865), .A2(new_n866), .B1(new_n424), .B2(new_n417), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n402), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n389), .A2(new_n866), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n405), .A2(new_n873), .A3(new_n869), .A4(new_n418), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n862), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n867), .ZN(new_n878));
  INV_X1    g0678(.A(new_n403), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n619), .A2(KEYINPUT72), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n405), .A2(new_n404), .A3(new_n406), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n882), .B2(new_n610), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n870), .A2(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n874), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n861), .B1(new_n877), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n405), .A2(new_n873), .A3(new_n418), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n874), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n873), .B1(new_n426), .B2(new_n620), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n862), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n887), .A2(new_n861), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n888), .A2(new_n894), .A3(KEYINPUT98), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT98), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n868), .A2(new_n862), .A3(new_n876), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n887), .A2(new_n893), .A3(new_n861), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n860), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n642), .A2(new_n653), .A3(new_n815), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n814), .B(KEYINPUT97), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n266), .A2(new_n653), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n305), .A2(new_n308), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n299), .B2(new_n304), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n897), .A2(new_n898), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n912), .A2(new_n913), .B1(new_n620), .B2(new_n866), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n731), .A2(new_n624), .A3(new_n723), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n623), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT99), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n700), .A2(new_n920), .A3(new_n678), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n705), .B1(KEYINPUT99), .B2(KEYINPUT31), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n715), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n817), .B1(new_n909), .B2(new_n910), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n897), .C2(new_n898), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT40), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n887), .A2(new_n893), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n929), .A2(new_n624), .A3(new_n923), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n624), .B2(new_n923), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n930), .A2(new_n931), .A3(new_n645), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n206), .B2(new_n736), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n919), .A2(new_n932), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n853), .B(new_n857), .C1(new_n934), .C2(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n749), .A2(new_n238), .ZN(new_n937));
  INV_X1    g0737(.A(new_n347), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n756), .B1(new_n671), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n740), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n744), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n599), .A2(new_n652), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n639), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n595), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n370), .B1(new_n768), .B2(new_n540), .ZN(new_n945));
  INV_X1    g0745(.A(G317), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n798), .A2(new_n771), .B1(new_n777), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(new_n785), .C2(G283), .ZN(new_n948));
  INV_X1    g0748(.A(G303), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n763), .A2(new_n949), .B1(new_n765), .B2(new_n789), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n761), .A2(new_n538), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G107), .B2(new_n775), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT108), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G159), .A2(new_n827), .B1(new_n769), .B2(new_n225), .ZN(new_n957));
  INV_X1    g0757(.A(G137), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n958), .B2(new_n777), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G50), .B2(new_n785), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n775), .A2(G68), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n765), .A2(new_n962), .B1(new_n761), .B2(new_n322), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n370), .B(new_n963), .C1(G150), .C2(new_n793), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n956), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n940), .B1(new_n941), .B2(new_n944), .C1(new_n967), .C2(new_n826), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n969));
  NAND3_X1  g0769(.A1(new_n625), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT100), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n531), .B2(new_n653), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n652), .B1(new_n529), .B2(new_n530), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n970), .A2(new_n972), .B1(new_n640), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n969), .B1(new_n669), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n667), .B1(new_n659), .B2(new_n661), .ZN(new_n977));
  INV_X1    g0777(.A(new_n969), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n977), .A2(new_n665), .A3(new_n974), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n669), .B2(new_n975), .ZN(new_n982));
  OAI211_X1 g0782(.A(KEYINPUT44), .B(new_n974), .C1(new_n977), .C2(new_n665), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n663), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT106), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT106), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n980), .A2(new_n984), .A3(new_n987), .A4(new_n663), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n715), .B1(new_n713), .B2(KEYINPUT88), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n709), .B(new_n691), .C1(new_n711), .C2(new_n712), .ZN(new_n991));
  OAI21_X1  g0791(.A(G330), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT105), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n730), .A2(KEYINPUT89), .ZN(new_n994));
  INV_X1    g0794(.A(new_n729), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n723), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n662), .A2(new_n668), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n656), .A2(new_n997), .A3(new_n977), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n656), .B1(new_n997), .B2(new_n977), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n992), .A2(new_n993), .A3(new_n996), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n980), .A2(new_n984), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n663), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n989), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n993), .B1(new_n732), .B2(new_n1000), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n732), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n672), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n738), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1003), .A2(new_n975), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT102), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n531), .B1(new_n974), .B2(new_n480), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n653), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n977), .A2(new_n975), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT101), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT103), .Z(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1013), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1029), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n1012), .A3(new_n1027), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n968), .B1(new_n1010), .B2(new_n1033), .ZN(G387));
  OR2_X1    g0834(.A1(new_n662), .A2(new_n941), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n746), .A2(new_n674), .B1(G107), .B2(new_n210), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n235), .A2(G45), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n674), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n1038), .C1(G68), .C2(G77), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n345), .A2(new_n202), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT50), .Z(new_n1041));
  AOI21_X1  g0841(.A(new_n750), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1036), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n739), .B1(new_n1043), .B2(new_n756), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT109), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G322), .A2(new_n791), .B1(new_n827), .B2(G311), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n946), .B2(new_n763), .C1(new_n784), .C2(new_n949), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT48), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT48), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n799), .A2(new_n794), .B1(G283), .B2(new_n775), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n768), .A2(new_n538), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n310), .B(new_n1056), .C1(G326), .C2(new_n796), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n778), .A2(new_n765), .B1(new_n781), .B2(new_n252), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n370), .B(new_n1059), .C1(G97), .C2(new_n769), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n763), .A2(new_n202), .B1(new_n777), .B2(new_n837), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n225), .B2(new_n794), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n582), .A2(new_n775), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n827), .A2(new_n327), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1045), .B1(new_n1066), .B2(new_n754), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1000), .A2(new_n738), .B1(new_n1035), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n732), .A2(new_n1000), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n672), .B(KEYINPUT110), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n732), .A2(new_n1000), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(G393));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1004), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1002), .A2(KEYINPUT111), .A3(new_n1003), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1075), .A2(new_n1076), .B1(new_n988), .B2(new_n986), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n974), .A2(new_n744), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n370), .B1(new_n768), .B2(new_n353), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G283), .A2(new_n794), .B1(new_n796), .B2(G322), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n430), .B2(new_n781), .C1(new_n949), .C2(new_n771), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(G116), .C2(new_n775), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n763), .A2(new_n789), .B1(new_n765), .B2(new_n946), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n763), .A2(new_n778), .B1(new_n765), .B2(new_n837), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n345), .B2(new_n785), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n370), .B(new_n830), .C1(G50), .C2(new_n827), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n261), .B2(new_n833), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n761), .A2(new_n252), .B1(new_n777), .B2(new_n962), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT112), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1082), .A2(new_n1084), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n826), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n749), .A2(new_n246), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n756), .B1(G97), .B2(new_n671), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n740), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1077), .A2(new_n738), .B1(new_n1078), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n732), .A2(new_n1000), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1070), .B1(new_n1077), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(G390));
  OAI211_X1 g0903(.A(G330), .B(new_n815), .C1(new_n990), .C2(new_n991), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n911), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n923), .A2(new_n924), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n645), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n811), .A2(new_n815), .A3(new_n911), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n728), .A2(new_n653), .A3(new_n815), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n905), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n816), .A2(G330), .A3(new_n923), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n1105), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1110), .A2(new_n906), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n923), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n624), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n623), .A2(new_n917), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT98), .B1(new_n888), .B2(new_n894), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n899), .A2(new_n896), .A3(new_n900), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n912), .A2(new_n859), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1113), .A2(new_n911), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n859), .B(KEYINPUT113), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n928), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1123), .A2(new_n1111), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1116), .A2(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1108), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n1111), .A3(new_n1126), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1119), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1115), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1108), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n906), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1129), .A2(new_n1070), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1120), .A2(new_n1121), .A3(new_n742), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n824), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n739), .B1(new_n327), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n793), .A2(G132), .B1(new_n769), .B2(G50), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n765), .C1(new_n958), .C2(new_n771), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n310), .B1(new_n777), .B2(new_n1147), .C1(new_n833), .C2(new_n778), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n761), .A2(new_n837), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT54), .B(G143), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1149), .B(new_n1151), .C1(new_n784), .C2(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n784), .A2(new_n540), .B1(new_n353), .B2(new_n771), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT114), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G68), .A2(new_n769), .B1(new_n796), .B2(G294), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n793), .A2(G116), .B1(new_n791), .B2(G283), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n833), .A2(new_n261), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1158), .A2(new_n310), .A3(new_n762), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1154), .A2(KEYINPUT114), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1153), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1143), .B1(new_n1162), .B2(new_n754), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1140), .A2(new_n738), .B1(new_n1141), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1139), .A2(new_n1164), .ZN(G378));
  AOI21_X1  g0965(.A(new_n740), .B1(new_n202), .B2(new_n824), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n796), .A2(G283), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n353), .B2(new_n763), .C1(new_n538), .C2(new_n765), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G41), .B(new_n310), .C1(new_n794), .C2(new_n225), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n827), .B1(new_n769), .B2(G58), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n961), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n781), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1169), .B(new_n1172), .C1(new_n582), .C2(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n202), .B1(new_n270), .B2(G41), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OR3_X1    g0978(.A1(new_n761), .A2(new_n1152), .A3(KEYINPUT115), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT115), .B1(new_n761), .B2(new_n1152), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n1145), .C2(new_n763), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT116), .Z(new_n1182));
  OAI22_X1  g0982(.A1(new_n1147), .A2(new_n765), .B1(new_n781), .B2(new_n958), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n833), .A2(new_n837), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G132), .C2(new_n827), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n778), .B2(new_n768), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1178), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n826), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT117), .Z(new_n1194));
  NAND3_X1  g0994(.A1(new_n342), .A2(new_n334), .A3(new_n866), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n334), .A2(new_n866), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n336), .B(new_n1196), .C1(new_n340), .C2(new_n341), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1167), .B(new_n1194), .C1(new_n1201), .C2(new_n742), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1201), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n929), .B2(G330), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1107), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n877), .A2(new_n887), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT40), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n619), .A2(new_n403), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n389), .B(new_n866), .C1(new_n1208), .C2(new_n610), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n890), .A2(new_n874), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT38), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n876), .B1(new_n427), .B2(new_n878), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(KEYINPUT38), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT40), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1207), .A2(new_n1215), .A3(new_n645), .A4(new_n1201), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n859), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1204), .A2(new_n1216), .B1(new_n1217), .B2(new_n914), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n925), .A2(new_n926), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n927), .A2(new_n928), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(G330), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1201), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n929), .A2(G330), .A3(new_n1203), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n902), .A3(new_n915), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1202), .B1(new_n1225), .B2(new_n738), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1138), .A2(new_n1133), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1070), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1138), .A2(new_n1133), .B1(new_n1224), .B2(new_n1218), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT57), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1229), .B2(new_n1231), .ZN(G375));
  OAI211_X1 g1032(.A(new_n1119), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT118), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1110), .A2(new_n906), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1119), .B1(new_n1237), .B2(new_n1134), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .A4(new_n1008), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n739), .B1(G68), .B2(new_n1142), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n763), .A2(new_n958), .B1(new_n771), .B2(new_n1152), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n370), .B(new_n1242), .C1(G58), .C2(new_n769), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1173), .A2(G150), .B1(new_n796), .B2(G128), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G132), .A2(new_n791), .B1(new_n794), .B2(G159), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n775), .A2(G50), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n793), .A2(G283), .B1(new_n827), .B2(G116), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n791), .A2(G294), .B1(new_n796), .B2(G303), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n540), .C2(new_n761), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n370), .B1(new_n768), .B2(new_n261), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT119), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1063), .C1(new_n353), .C2(new_n784), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1241), .B1(new_n1254), .B2(new_n754), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT120), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n911), .B2(new_n743), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1116), .B2(new_n737), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1240), .A2(new_n1258), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT121), .Z(G381));
  INV_X1    g1060(.A(new_n1226), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1070), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1230), .B2(KEYINPUT57), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1119), .B1(new_n1140), .B2(new_n1137), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1218), .A2(new_n1224), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1261), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1271));
  OR4_X1    g1071(.A1(G387), .A2(G381), .A3(new_n1270), .A4(new_n1271), .ZN(G407));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  OAI211_X1 g1073(.A(G390), .B(new_n968), .C1(new_n1010), .C2(new_n1033), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT124), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n807), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1274), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1275), .A2(new_n1279), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT125), .ZN(new_n1285));
  INV_X1    g1085(.A(G213), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(G343), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1237), .A2(KEYINPUT118), .A3(new_n1119), .A4(new_n1134), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1235), .B(new_n1290), .C1(new_n1238), .C2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT122), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1116), .A2(new_n1293), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1119), .A4(new_n1134), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1262), .B1(new_n1295), .B2(KEYINPUT122), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1258), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(G384), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G384), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(KEYINPUT123), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1291), .B1(new_n1137), .B2(new_n1133), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1236), .A2(new_n1302), .A3(new_n1239), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT122), .B1(new_n1233), .B2(new_n1291), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(new_n1070), .A3(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1298), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(KEYINPUT123), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1289), .B1(new_n1301), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT123), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1305), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1258), .B1(new_n1312), .B2(new_n1292), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1313), .B2(G384), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1314), .A2(new_n1288), .A3(new_n1308), .A4(new_n1299), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1139), .A2(new_n1164), .A3(new_n1226), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1230), .A2(new_n1009), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1287), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1310), .A2(new_n1315), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1314), .A2(new_n1308), .A3(new_n1299), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1287), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1139), .A2(new_n1226), .A3(new_n1164), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1265), .A2(new_n1008), .A3(new_n1266), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(G375), .B2(G378), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT123), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1299), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1328), .A2(new_n1331), .A3(KEYINPUT63), .A4(new_n1308), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1285), .A2(new_n1320), .A3(new_n1323), .A4(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT62), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1328), .A2(new_n1331), .A3(new_n1336), .A4(new_n1308), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1335), .A2(new_n1282), .A3(new_n1337), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1310), .A2(new_n1315), .A3(new_n1319), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1334), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1333), .A2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(KEYINPUT126), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1283), .B(new_n1281), .C1(new_n1322), .C2(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1334), .A2(KEYINPUT126), .A3(new_n1308), .A4(new_n1331), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1268), .B(G378), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1345), .B(new_n1346), .ZN(G402));
endmodule


