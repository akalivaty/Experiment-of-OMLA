//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n457), .B1(new_n448), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(KEYINPUT3), .A3(new_n469), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n461), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NOR2_X1   g060(.A1(new_n473), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  OR3_X1    g063(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n472), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n461), .A2(new_n463), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR4_X1   g070(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n495), .A4(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n472), .A2(new_n461), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n498), .A2(KEYINPUT68), .A3(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT69), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n506), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(new_n504), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n509), .A2(new_n514), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n513), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(new_n523), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n504), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(G90), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  XOR2_X1   g111(.A(KEYINPUT71), .B(G81), .Z(new_n537));
  NAND2_X1  g112(.A1(new_n513), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n508), .A2(G43), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n504), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n513), .A2(G91), .B1(G651), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n508), .A2(G53), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G299));
  NAND2_X1  g135(.A1(new_n508), .A2(G49), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n513), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  AND2_X1   g139(.A1(G48), .A2(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n506), .A2(new_n507), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n551), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n566), .A2(KEYINPUT73), .B1(new_n569), .B2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n513), .A2(G86), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n506), .A2(new_n572), .A3(new_n507), .A4(new_n565), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(G47), .A2(new_n508), .B1(new_n513), .B2(G85), .ZN(new_n575));
  NAND2_X1  g150(.A1(G72), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G60), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n551), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n504), .B1(new_n578), .B2(KEYINPUT74), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(KEYINPUT74), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(new_n513), .A2(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n551), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n508), .A2(G54), .B1(G651), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G171), .B2(new_n592), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(G171), .B2(new_n592), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n559), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(new_n559), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(new_n591), .ZN(new_n599));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g180(.A(new_n494), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n470), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n478), .A2(G135), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n480), .A2(G123), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT75), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n613), .A2(new_n473), .A3(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n473), .B2(G111), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n611), .B(new_n612), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n630), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT77), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT17), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n641), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n639), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n641), .A3(new_n637), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  INV_X1    g223(.A(new_n641), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(new_n637), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n646), .B(new_n648), .C1(new_n640), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT20), .Z(new_n662));
  OR2_X1    g237(.A1(new_n655), .A2(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n660), .A3(new_n658), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n660), .C2(new_n663), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G27), .A2(G29), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(G164), .B2(G29), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(G2078), .ZN(new_n674));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G35), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G162), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT29), .Z(new_n678));
  INV_X1    g253(.A(G2090), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NOR2_X1   g256(.A1(G171), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(G5), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G1961), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n674), .B(new_n685), .C1(new_n684), .C2(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n675), .A2(G32), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n478), .A2(G141), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n480), .A2(G129), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT85), .B(KEYINPUT26), .Z(new_n690));
  NAND3_X1  g265(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n470), .A2(G105), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n688), .A2(new_n689), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n687), .B1(new_n695), .B2(new_n675), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT27), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1996), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n681), .A2(G19), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n543), .B2(new_n681), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1341), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n673), .A2(G2078), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n675), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT25), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n606), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n473), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G139), .B2(new_n478), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(new_n675), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G2072), .Z(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AOI21_X1  g286(.A(G29), .B1(new_n711), .B2(KEYINPUT24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(KEYINPUT24), .B2(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n475), .B2(new_n675), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2084), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n701), .A2(new_n702), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G28), .ZN(new_n717));
  OR2_X1    g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  NAND2_X1  g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n717), .A2(new_n675), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n617), .B2(new_n675), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT87), .Z(new_n722));
  NOR2_X1   g297(.A1(G4), .A2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n599), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G1348), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n681), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n681), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT86), .B(G1966), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G1348), .B2(new_n724), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n716), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT88), .B(KEYINPUT23), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n681), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G299), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1956), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n678), .A2(new_n679), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n675), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n478), .A2(G140), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT83), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G128), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT84), .B1(G104), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(KEYINPUT84), .A2(G104), .A3(G2105), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G116), .B2(new_n473), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n742), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n739), .A2(new_n740), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n686), .A2(new_n698), .A3(new_n733), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n681), .A2(G23), .ZN(new_n757));
  INV_X1    g332(.A(G288), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n681), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT82), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT33), .B(G1976), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n681), .A2(G22), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G166), .B2(new_n681), .ZN(new_n764));
  INV_X1    g339(.A(G1971), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G6), .B(G305), .S(G16), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT32), .B(G1981), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n762), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(KEYINPUT34), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n480), .A2(G119), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n473), .A2(G107), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G131), .B2(new_n478), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT80), .ZN(new_n778));
  MUX2_X1   g353(.A(G25), .B(new_n778), .S(G29), .Z(new_n779));
  XOR2_X1   g354(.A(KEYINPUT35), .B(G1991), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G24), .ZN(new_n782));
  XOR2_X1   g357(.A(G290), .B(KEYINPUT81), .Z(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n771), .A2(new_n772), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT36), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT36), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n756), .B1(new_n788), .B2(new_n789), .ZN(G311));
  INV_X1    g365(.A(G311), .ZN(G150));
  XNOR2_X1  g366(.A(KEYINPUT89), .B(G55), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n508), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n513), .A2(G93), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(new_n504), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT91), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT91), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G860), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT37), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n599), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n798), .A2(new_n542), .A3(new_n800), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n807));
  INV_X1    g382(.A(new_n797), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n542), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n543), .A2(KEYINPUT90), .A3(new_n797), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n805), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  INV_X1    g390(.A(G860), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(KEYINPUT39), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n803), .B1(new_n815), .B2(new_n817), .ZN(G145));
  XNOR2_X1  g393(.A(new_n617), .B(new_n475), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n484), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n822));
  AOI211_X1 g397(.A(new_n822), .B(new_n493), .C1(new_n501), .C2(new_n502), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n499), .A2(new_n500), .ZN(new_n824));
  INV_X1    g399(.A(new_n496), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n502), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n493), .ZN(new_n827));
  AOI21_X1  g402(.A(KEYINPUT92), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n751), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n695), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n827), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n822), .ZN(new_n833));
  NAND2_X1  g408(.A1(G164), .A2(KEYINPUT92), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n751), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n694), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n831), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n480), .A2(G130), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n473), .A2(G118), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G142), .B2(new_n478), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(new_n608), .Z(new_n845));
  OR2_X1    g420(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n778), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n839), .A2(new_n845), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n846), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n821), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n820), .A3(new_n850), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n859));
  NAND2_X1  g434(.A1(G299), .A2(new_n599), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n559), .A2(new_n591), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(KEYINPUT94), .A3(new_n861), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n559), .A2(new_n591), .A3(KEYINPUT94), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(KEYINPUT41), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n811), .B(new_n602), .Z(new_n869));
  OR2_X1    g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n866), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(G303), .B(G288), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT42), .Z(new_n882));
  NAND3_X1  g457(.A1(new_n875), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n876), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n870), .A3(new_n874), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n882), .A2(new_n876), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n859), .B(G868), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n883), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT97), .B1(new_n889), .B2(new_n592), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n801), .A2(new_n592), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G295));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G331));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  NAND2_X1  g469(.A1(G301), .A2(G286), .ZN(new_n895));
  OAI211_X1 g470(.A(G168), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n812), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n811), .A2(new_n895), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(new_n871), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(KEYINPUT99), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n811), .A2(new_n903), .A3(new_n895), .A4(new_n896), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n812), .A2(new_n897), .A3(KEYINPUT98), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT98), .B1(new_n812), .B2(new_n897), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n902), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n901), .B1(new_n907), .B2(new_n868), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n908), .B2(new_n881), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n871), .A2(new_n863), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n910), .B(new_n900), .C1(new_n863), .C2(new_n862), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n873), .B2(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n881), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n864), .A2(new_n867), .ZN(new_n918));
  INV_X1    g493(.A(new_n906), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n812), .A2(new_n897), .A3(KEYINPUT98), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n902), .A2(new_n904), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n914), .B1(new_n923), .B2(new_n901), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n916), .B1(new_n909), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT101), .B(new_n916), .C1(new_n909), .C2(new_n924), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n894), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n909), .A2(new_n915), .A3(KEYINPUT43), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n909), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(G397));
  NOR3_X1   g508(.A1(new_n823), .A2(new_n828), .A3(G1384), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n466), .A2(G2105), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n470), .A2(G101), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(G40), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n936), .A2(new_n474), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT103), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT104), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n935), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n785), .B1(new_n575), .B2(new_n580), .ZN(new_n946));
  NOR2_X1   g521(.A1(G290), .A2(G1986), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT105), .Z(new_n949));
  XNOR2_X1  g524(.A(new_n751), .B(new_n753), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n945), .A2(KEYINPUT107), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n950), .B(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n942), .A2(new_n944), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n694), .B(G1996), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n953), .A2(new_n957), .B1(new_n945), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n778), .B(new_n780), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n945), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n949), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1384), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n823), .A2(new_n828), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n826), .B2(new_n827), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n940), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n765), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n832), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n679), .A4(new_n940), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n964), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G303), .A2(G8), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n502), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT68), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(new_n496), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n973), .B1(new_n984), .B2(new_n493), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n939), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n964), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n566), .A2(KEYINPUT73), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n569), .A2(G651), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT109), .B(G86), .Z(new_n992));
  NAND4_X1  g567(.A1(new_n506), .A2(new_n507), .A3(new_n512), .A4(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n573), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G1981), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n570), .A2(new_n571), .A3(new_n996), .A4(new_n573), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(KEYINPUT49), .A3(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n989), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n758), .A2(G1976), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n989), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n940), .A2(new_n969), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n997), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G288), .A2(G1976), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1005), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n989), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n981), .A2(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n987), .B1(new_n985), .B2(new_n965), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n833), .A2(new_n834), .A3(new_n966), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1971), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n976), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n971), .A2(KEYINPUT112), .A3(new_n976), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n979), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT113), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1013), .B1(new_n980), .B2(new_n977), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(new_n979), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2078), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1021), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(G2078), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1021), .B(new_n1038), .C1(G164), .C2(new_n967), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n974), .A2(new_n975), .A3(new_n940), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n684), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G171), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(KEYINPUT120), .A3(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G164), .A2(new_n967), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n730), .B1(new_n970), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G2084), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n974), .A2(new_n975), .A3(new_n1050), .A4(new_n940), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(G168), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(G168), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1047), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1033), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT123), .B1(new_n1062), .B2(KEYINPUT62), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1064), .B(new_n1056), .C1(new_n1055), .C2(new_n1058), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1019), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1070), .A2(new_n1038), .A3(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1022), .B(new_n1072), .C1(new_n934), .C2(KEYINPUT45), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1037), .A2(new_n1073), .A3(new_n1041), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1037), .A2(new_n1039), .A3(G301), .A4(new_n1041), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(KEYINPUT54), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1062), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1031), .B1(new_n1027), .B2(new_n979), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n1082));
  NAND2_X1  g657(.A1(new_n557), .A2(new_n558), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n555), .A2(KEYINPUT116), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n555), .A2(KEYINPUT116), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n559), .A2(KEYINPUT57), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1040), .A2(new_n738), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1021), .A2(new_n1022), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1040), .A2(new_n726), .B1(new_n988), .B2(new_n753), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n591), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1088), .A3(new_n1087), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g675(.A(G1996), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1021), .A2(new_n1022), .A3(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1010), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n542), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1105), .B2(KEYINPUT118), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1098), .A2(new_n1093), .A3(new_n1109), .A4(KEYINPUT61), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1100), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT59), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1108), .B(new_n1110), .C1(new_n1106), .C2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1094), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1098), .A2(new_n1093), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1098), .B2(KEYINPUT119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1099), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1074), .A2(G171), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1045), .A2(new_n1046), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1081), .B(new_n1122), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1067), .A2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n964), .B(G286), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n977), .A2(new_n980), .ZN(new_n1137));
  AND4_X1   g712(.A1(KEYINPUT63), .A2(new_n1030), .A3(new_n1131), .A4(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n963), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n945), .A2(new_n1141), .A3(new_n947), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n942), .A2(new_n944), .A3(new_n947), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT48), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(KEYINPUT48), .A3(new_n1144), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n959), .A3(new_n962), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n780), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n778), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n744), .A2(new_n750), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n959), .A2(new_n1151), .B1(new_n753), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1153), .B2(new_n956), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n942), .A2(KEYINPUT46), .A3(new_n1101), .A4(new_n944), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT124), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n955), .A2(new_n695), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n942), .A2(new_n1101), .A3(new_n944), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1157), .A2(new_n945), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT125), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1156), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT47), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT47), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1162), .A2(new_n1167), .A3(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1154), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1140), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g745(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n857), .B(new_n1172), .C1(new_n927), .C2(new_n928), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


