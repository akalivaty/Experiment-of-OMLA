//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G116), .B2(G270), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G58), .A2(G232), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G50), .A2(G226), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n220), .A2(new_n223), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT65), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT64), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G107), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n247), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT69), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n253), .A2(new_n256), .A3(G1), .A4(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT66), .B(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(new_n261), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(G45), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(KEYINPUT67), .A3(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n254), .A2(G274), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n254), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G244), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n259), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G20), .A2(G77), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT15), .B(G87), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n226), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n278), .B1(new_n279), .B2(new_n280), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n227), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n285), .B(new_n227), .C1(G1), .C2(new_n226), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G77), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G77), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n276), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n277), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT12), .B1(new_n292), .B2(G68), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n289), .B2(G68), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n280), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n304), .A2(new_n305), .A3(new_n286), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n304), .B2(new_n286), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(KEYINPUT73), .B(new_n301), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  INV_X1    g0113(.A(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n248), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G232), .B2(new_n248), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n313), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n258), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n274), .A2(G238), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n272), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n272), .A2(new_n323), .A3(new_n327), .A4(new_n324), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(G190), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n312), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n328), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n326), .B2(new_n328), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n336), .B(new_n333), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n330), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n331), .A2(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n331), .A2(new_n346), .A3(G169), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n345), .B(new_n347), .C1(new_n348), .C2(new_n331), .ZN(new_n349));
  INV_X1    g0149(.A(new_n312), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G222), .A2(G1698), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n248), .A2(G223), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n247), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n321), .A2(new_n303), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT68), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n258), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n274), .A2(G226), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n272), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n296), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n203), .A2(G20), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  INV_X1    g0165(.A(G58), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT70), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G58), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT8), .ZN(new_n370));
  OR2_X1    g0170(.A1(KEYINPUT8), .A2(G58), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n364), .B1(new_n365), .B2(new_n282), .C1(new_n372), .C2(new_n280), .ZN(new_n373));
  INV_X1    g0173(.A(new_n292), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n286), .B1(new_n202), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n289), .A2(G50), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n363), .B(new_n377), .C1(G179), .C2(new_n362), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n343), .A2(new_n351), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n362), .A2(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(KEYINPUT9), .A3(new_n376), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n360), .A2(G190), .A3(new_n272), .A4(new_n361), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT10), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n375), .A2(KEYINPUT9), .A3(new_n376), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT9), .B1(new_n375), .B2(new_n376), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT10), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n382), .A4(new_n384), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n298), .B(new_n379), .C1(new_n386), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n247), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n216), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n282), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT70), .B(G58), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n201), .B1(new_n402), .B2(G68), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(new_n226), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n394), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n321), .B2(new_n226), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n395), .B(G20), .C1(new_n318), .C2(new_n320), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n367), .A2(new_n369), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n224), .B1(new_n409), .B2(new_n216), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n400), .B1(new_n410), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n412), .A3(new_n286), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT75), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n370), .A2(new_n288), .A3(new_n371), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n374), .B1(new_n370), .B2(new_n371), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n372), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n415), .B(KEYINPUT75), .C1(new_n419), .C2(new_n374), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n274), .A2(G232), .ZN(new_n423));
  OR2_X1    g0223(.A1(G223), .A2(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n314), .A2(G1698), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n318), .A2(new_n424), .A3(new_n320), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n258), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n272), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n335), .ZN(new_n431));
  INV_X1    g0231(.A(G190), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n272), .A2(new_n429), .A3(new_n432), .A4(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n393), .B1(new_n422), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n413), .A3(new_n421), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(G169), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n272), .A2(new_n429), .A3(G179), .A4(new_n423), .ZN(new_n441));
  AOI221_X4 g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .C1(new_n413), .C2(new_n421), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n413), .A2(new_n421), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT18), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n438), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n276), .A2(G200), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n259), .A2(G190), .A3(new_n272), .A4(new_n275), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n291), .A4(new_n294), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n265), .A2(new_n267), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n261), .B(G45), .C1(new_n455), .C2(G41), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(new_n254), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n262), .A2(new_n455), .ZN(new_n459));
  INV_X1    g0259(.A(new_n457), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(G274), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT76), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(new_n248), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n258), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT76), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n458), .A2(new_n461), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n463), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n476), .A2(new_n477), .A3(G107), .ZN(new_n478));
  XNOR2_X1  g0278(.A(G97), .B(G107), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n480), .A2(new_n226), .B1(new_n303), .B2(new_n282), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n251), .B1(new_n396), .B2(new_n397), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n286), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n286), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n261), .A2(G33), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n292), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n292), .A2(G97), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n483), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n462), .B1(new_n258), .B2(new_n470), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n475), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n471), .A2(new_n461), .A3(new_n458), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n296), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n463), .A2(new_n348), .A3(new_n471), .A4(new_n473), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(new_n488), .A3(new_n490), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n217), .A2(new_n248), .ZN(new_n501));
  INV_X1    g0301(.A(G244), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n318), .A2(new_n501), .A3(new_n320), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT78), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n255), .A2(new_n257), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n269), .A2(KEYINPUT77), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n269), .A2(KEYINPUT77), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(G250), .A3(new_n254), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n261), .A2(G45), .A3(G274), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n296), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n280), .B2(new_n477), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n247), .A2(new_n226), .A3(G68), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n517), .C1(new_n280), .C2(new_n477), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n226), .B1(new_n313), .B2(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n208), .A2(new_n477), .A3(new_n251), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n519), .A2(new_n520), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n286), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n279), .A2(new_n374), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n279), .C2(new_n486), .ZN(new_n529));
  INV_X1    g0329(.A(new_n508), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n258), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n515), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n516), .B(new_n529), .C1(G179), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n487), .A2(G87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n528), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(G200), .B1(new_n510), .B2(new_n515), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(G190), .A3(new_n533), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n500), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n318), .A2(new_n320), .A3(new_n226), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n247), .A2(new_n547), .A3(new_n226), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n226), .A2(G107), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT23), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n549), .A2(KEYINPUT24), .A3(new_n550), .A4(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n286), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n486), .A2(new_n251), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n247), .A2(G257), .A3(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G294), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n318), .A2(new_n320), .A3(G250), .A4(new_n248), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n258), .ZN(new_n565));
  OAI211_X1 g0365(.A(G264), .B(new_n254), .C1(new_n456), .C2(new_n457), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n461), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n335), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(KEYINPUT81), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n461), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(new_n572), .A3(new_n258), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n568), .B1(new_n574), .B2(G190), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT80), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(KEYINPUT25), .C1(new_n292), .C2(G107), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n576), .A2(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(KEYINPUT25), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n374), .A2(new_n578), .A3(new_n251), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n560), .A2(new_n575), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n571), .A2(G179), .A3(new_n565), .ZN(new_n582));
  INV_X1    g0382(.A(new_n573), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n572), .B1(new_n564), .B2(new_n258), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n583), .A2(new_n570), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n582), .B1(new_n585), .B2(new_n296), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n557), .A2(new_n577), .A3(new_n559), .A4(new_n580), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n374), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n484), .A2(G116), .A3(new_n292), .A4(new_n485), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n285), .A2(new_n227), .B1(G20), .B2(new_n589), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n468), .B(new_n226), .C1(G33), .C2(new_n477), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n590), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n318), .A2(new_n320), .A3(G257), .A4(new_n248), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n318), .A2(new_n320), .A3(G264), .A4(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n247), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n258), .ZN(new_n601));
  OAI211_X1 g0401(.A(G270), .B(new_n254), .C1(new_n456), .C2(new_n457), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n461), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n596), .B(G169), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(new_n258), .ZN(new_n607));
  AND4_X1   g0407(.A1(G179), .A2(new_n607), .A3(new_n461), .A4(new_n602), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n596), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n461), .A3(new_n602), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(KEYINPUT21), .A3(G169), .A4(new_n596), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n596), .B1(new_n610), .B2(G200), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n432), .B2(new_n610), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n588), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n544), .A2(new_n581), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n392), .A2(new_n454), .A3(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n343), .A2(new_n298), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n438), .B1(new_n618), .B2(new_n351), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n391), .A2(new_n386), .A3(KEYINPUT82), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT82), .B1(new_n391), .B2(new_n386), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n619), .A2(new_n449), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n378), .ZN(new_n623));
  INV_X1    g0423(.A(new_n535), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n542), .B2(new_n499), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(KEYINPUT26), .A3(new_n535), .A4(new_n541), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n588), .A2(new_n612), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n500), .A3(new_n581), .A4(new_n543), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n392), .A2(new_n454), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(G369));
  NAND2_X1  g0434(.A1(new_n612), .A2(new_n614), .ZN(new_n635));
  INV_X1    g0435(.A(G13), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n261), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n640), .A3(new_n261), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n639), .A2(G213), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G343), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n596), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n612), .A2(new_n596), .A3(new_n644), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(G330), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n612), .A2(new_n644), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n587), .B1(new_n586), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n581), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n586), .A2(new_n587), .A3(new_n644), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n644), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n586), .A2(new_n587), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n649), .A2(new_n581), .A3(new_n651), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n221), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n262), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n524), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n225), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  INV_X1    g0466(.A(new_n610), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n458), .A2(new_n461), .A3(new_n472), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n472), .B1(new_n458), .B2(new_n461), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n670), .B2(new_n471), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n348), .A3(new_n567), .A4(new_n534), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT84), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(KEYINPUT84), .A2(KEYINPUT30), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n608), .A2(new_n565), .A3(new_n566), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n492), .A2(new_n533), .A3(new_n532), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n565), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n610), .A2(new_n682), .A3(new_n348), .A4(new_n677), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n495), .A2(new_n534), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n566), .A4(new_n675), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n672), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT31), .B1(new_n686), .B2(new_n644), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT85), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n644), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT85), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n544), .A2(new_n581), .A3(new_n615), .A4(new_n656), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n632), .A2(new_n656), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n644), .B1(new_n629), .B2(new_n631), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n666), .B1(new_n706), .B2(G1), .ZN(G364));
  NAND2_X1  g0507(.A1(new_n637), .A2(G45), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n662), .A2(G1), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT87), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT87), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n646), .A2(new_n647), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n717), .B2(KEYINPUT86), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n648), .B1(new_n717), .B2(KEYINPUT86), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n713), .B(KEYINPUT88), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n660), .A2(new_n247), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n240), .B2(G45), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G45), .B2(new_n225), .ZN(new_n726));
  INV_X1    g0526(.A(G355), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n247), .A2(new_n221), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n726), .B1(G116), .B2(new_n221), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n636), .A2(new_n317), .A3(KEYINPUT89), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT89), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G13), .B2(G33), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n227), .B1(G20), .B2(new_n296), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n736), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n226), .A2(new_n432), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n335), .A2(G179), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(KEYINPUT91), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(KEYINPUT91), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n226), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n749), .A2(G303), .B1(G329), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n226), .B1(new_n751), .B2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G294), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n348), .A2(new_n335), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n758), .A2(new_n750), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n348), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n740), .A2(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT92), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n741), .A2(new_n750), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n750), .A2(new_n763), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n321), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n740), .A2(new_n758), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n769), .B(new_n772), .C1(G326), .C2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n754), .A2(new_n757), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT32), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n753), .B2(G159), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n760), .A2(new_n216), .B1(new_n409), .B2(new_n764), .ZN(new_n778));
  INV_X1    g0578(.A(new_n770), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n777), .B(new_n778), .C1(G77), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n767), .A2(new_n251), .ZN(new_n781));
  INV_X1    g0581(.A(new_n773), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n247), .B1(new_n782), .B2(new_n202), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n781), .B(new_n783), .C1(G97), .C2(new_n756), .ZN(new_n784));
  INV_X1    g0584(.A(new_n745), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n753), .A2(new_n776), .A3(G159), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n780), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n739), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n738), .B(new_n789), .C1(new_n714), .C2(new_n735), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n719), .A2(new_n720), .B1(new_n722), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  AND2_X1   g0592(.A1(new_n295), .A2(new_n297), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n644), .A2(new_n295), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(new_n277), .B1(new_n453), .B2(new_n794), .ZN(new_n795));
  AND4_X1   g0595(.A1(new_n295), .A2(new_n656), .A3(new_n297), .A4(new_n277), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT93), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT93), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n793), .A2(new_n277), .A3(new_n656), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n453), .A2(new_n794), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n298), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n699), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n797), .A2(new_n801), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n632), .A2(new_n656), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n698), .B(new_n806), .Z(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n713), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n721), .B1(new_n802), .B2(new_n733), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n733), .A2(new_n736), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n303), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n247), .B1(new_n749), .B2(G107), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n773), .A2(G303), .B1(new_n756), .B2(G97), .ZN(new_n813));
  INV_X1    g0613(.A(new_n767), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G87), .A2(new_n814), .B1(new_n753), .B2(G311), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n779), .A2(G116), .B1(new_n759), .B2(G283), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n764), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G294), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G143), .A2(new_n818), .B1(new_n779), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n823), .B2(new_n782), .C1(new_n365), .C2(new_n760), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT34), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n820), .B1(new_n821), .B2(new_n752), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n321), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n748), .B2(new_n202), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n402), .C2(new_n756), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n736), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n809), .A2(new_n811), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n808), .A2(new_n831), .ZN(G384));
  NAND2_X1  g0632(.A1(new_n805), .A2(new_n799), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n343), .B(new_n351), .C1(new_n312), .C2(new_n656), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT74), .B1(new_n341), .B2(new_n330), .ZN(new_n835));
  AND4_X1   g0635(.A1(KEYINPUT74), .A2(new_n330), .A3(new_n334), .A4(new_n337), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n351), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n656), .A2(new_n312), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n435), .A2(new_n437), .B1(new_n442), .B2(new_n446), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n415), .B1(new_n419), .B2(new_n374), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n413), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n642), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n445), .B2(new_n642), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n436), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n413), .A2(new_n421), .B1(new_n440), .B2(new_n441), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT94), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n444), .A2(new_n445), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT94), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT95), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n444), .B2(new_n642), .ZN(new_n856));
  INV_X1    g0656(.A(new_n642), .ZN(new_n857));
  AOI211_X1 g0657(.A(KEYINPUT95), .B(new_n857), .C1(new_n413), .C2(new_n421), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n436), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n848), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n845), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n845), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n841), .A2(new_n863), .B1(new_n448), .B2(new_n642), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT96), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT39), .B1(new_n861), .B2(new_n862), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n845), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n436), .A2(KEYINPUT97), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT97), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n434), .A2(new_n870), .A3(new_n413), .A4(new_n421), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n852), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n856), .A2(new_n858), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n444), .A2(new_n642), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT95), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n444), .A2(new_n855), .A3(new_n642), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(new_n436), .A3(new_n853), .A4(new_n851), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n874), .A2(new_n879), .B1(new_n842), .B2(new_n873), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n867), .B(new_n868), .C1(new_n880), .C2(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n866), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n349), .A2(new_n350), .A3(new_n656), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n864), .A2(KEYINPUT96), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n865), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n687), .A2(new_n688), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n802), .B1(new_n889), .B2(new_n696), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n840), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n867), .B1(new_n880), .B2(KEYINPUT38), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(KEYINPUT40), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n890), .B(new_n840), .C1(new_n862), .C2(new_n861), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n891), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n889), .A2(new_n696), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n454), .A3(new_n392), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n891), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n894), .A2(new_n895), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(G330), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n392), .A2(G330), .A3(new_n454), .A4(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n888), .B(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n392), .A2(new_n701), .A3(new_n454), .A4(new_n703), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n623), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n261), .B2(new_n637), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n226), .B(new_n227), .C1(new_n480), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(G116), .C1(new_n910), .C2(new_n480), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n303), .B(new_n225), .C1(new_n402), .C2(G68), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n216), .A2(G50), .ZN(new_n915));
  OAI211_X1 g0715(.A(G1), .B(new_n636), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT99), .ZN(G367));
  NAND2_X1  g0718(.A1(new_n708), .A2(G1), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n652), .A2(new_n653), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n650), .C1(new_n715), .C2(new_n714), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n922), .A2(new_n655), .A3(new_n658), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n698), .A2(new_n704), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n644), .A2(new_n498), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n494), .A2(new_n499), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n627), .A2(new_n644), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n658), .A2(new_n657), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n658), .A2(KEYINPUT45), .A3(new_n657), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n936), .B(new_n929), .C1(new_n658), .C2(new_n657), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n658), .A2(new_n657), .ZN(new_n939));
  INV_X1    g0739(.A(new_n929), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  AND4_X1   g0742(.A1(new_n655), .A2(new_n934), .A3(new_n938), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n937), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n655), .B1(new_n945), .B2(new_n934), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT104), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n698), .A2(new_n704), .A3(new_n923), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n925), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n925), .A2(new_n947), .A3(KEYINPUT105), .A4(new_n949), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n705), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n661), .B(KEYINPUT41), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n920), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n644), .A2(new_n537), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT100), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(new_n542), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n499), .B1(new_n927), .B2(new_n588), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(new_n656), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT42), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n658), .A2(new_n964), .A3(new_n927), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n658), .B2(new_n927), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n961), .B(KEYINPUT102), .C1(new_n963), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT102), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n960), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n970), .A3(new_n960), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT101), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT101), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n968), .A2(new_n973), .A3(new_n977), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n655), .A2(new_n940), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n957), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n785), .A2(new_n402), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n773), .A2(G143), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n756), .A2(G68), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n818), .A2(G150), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n779), .A2(G50), .B1(new_n759), .B2(G159), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT106), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n247), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n767), .A2(new_n303), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n752), .A2(new_n823), .ZN(new_n992));
  NOR4_X1   g0792(.A1(new_n987), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n782), .A2(new_n771), .B1(new_n477), .B2(new_n767), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT46), .B1(new_n748), .B2(new_n589), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n589), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n247), .B1(new_n759), .B2(G294), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n818), .A2(G303), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n753), .A2(G317), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n994), .B(new_n1001), .C1(G107), .C2(new_n756), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n779), .A2(G283), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n993), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT47), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n736), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n721), .B1(new_n960), .B2(new_n735), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n737), .B1(new_n221), .B2(new_n279), .C1(new_n236), .C2(new_n724), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n982), .A2(new_n1009), .ZN(G387));
  AOI22_X1  g0810(.A1(G322), .A2(new_n773), .B1(new_n759), .B2(G311), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n818), .A2(G317), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n599), .C2(new_n770), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1014));
  INV_X1    g0814(.A(G294), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n768), .B2(new_n755), .C1(new_n1015), .C2(new_n745), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT49), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n247), .B1(new_n753), .B2(G326), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n589), .C2(new_n767), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n785), .A2(G77), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n782), .A2(new_n399), .B1(new_n760), .B2(new_n372), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n818), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n365), .C2(new_n752), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n755), .A2(new_n279), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n247), .B1(new_n770), .B2(new_n216), .C1(new_n477), .C2(new_n767), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n739), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(G45), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n723), .B1(new_n233), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n663), .B2(new_n728), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n283), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n663), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n660), .A2(new_n251), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n735), .B(new_n736), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1027), .A2(new_n721), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n921), .A2(new_n735), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1038), .A2(new_n1039), .B1(new_n919), .B2(new_n923), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n661), .B1(new_n706), .B2(new_n923), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n924), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  NAND2_X1  g0843(.A1(new_n952), .A2(new_n953), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n947), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n924), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n661), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n947), .A2(new_n919), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n245), .A2(new_n723), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1049), .B(new_n737), .C1(new_n477), .C2(new_n221), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT107), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n818), .A2(G311), .B1(new_n773), .B2(G317), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT108), .B(KEYINPUT52), .Z(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n781), .B(new_n1054), .C1(G294), .C2(new_n779), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n753), .A2(G322), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n247), .B1(new_n759), .B2(G303), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n785), .A2(G283), .B1(G116), .B2(new_n756), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n782), .A2(new_n365), .B1(new_n764), .B2(new_n399), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n321), .B1(new_n785), .B2(G68), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G87), .A2(new_n814), .B1(new_n753), .B2(G143), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n755), .A2(new_n303), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n770), .A2(new_n283), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G50), .C2(new_n759), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1051), .B1(new_n1068), .B2(new_n736), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n940), .A2(new_n735), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1050), .A2(KEYINPUT107), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n722), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1047), .A2(new_n1048), .A3(new_n1072), .ZN(G390));
  NAND3_X1  g0873(.A1(new_n866), .A2(KEYINPUT109), .A3(new_n881), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n892), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n884), .B1(new_n833), .B2(new_n840), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n834), .A2(new_n839), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n796), .B1(new_n702), .B2(new_n804), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n883), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT109), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n866), .A2(new_n1081), .A3(new_n881), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT110), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n890), .A2(G330), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1078), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT110), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1077), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n799), .A2(new_n805), .B1(new_n834), .B2(new_n839), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1091), .A2(new_n892), .A3(new_n884), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1092), .A2(new_n1074), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n697), .A2(G330), .A3(new_n804), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n1078), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT111), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT111), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1095), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1084), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1090), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n906), .A2(new_n902), .A3(new_n623), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1094), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n841), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n841), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1086), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1105), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1090), .A2(new_n1096), .A3(new_n1099), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n661), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n745), .A2(new_n365), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n753), .A2(G125), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n767), .A2(new_n202), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n247), .B1(new_n755), .B2(new_n399), .C1(new_n782), .C2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT112), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1117), .B(new_n1119), .C1(new_n779), .C2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G132), .A2(new_n818), .B1(new_n759), .B2(G137), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1115), .A2(new_n1116), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n782), .A2(new_n768), .B1(new_n764), .B2(new_n589), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n321), .B1(new_n748), .B2(new_n208), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT113), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G294), .C2(new_n753), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n759), .A2(G107), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n779), .A2(G97), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1128), .A2(new_n820), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1124), .B1(new_n1131), .B2(new_n1064), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n736), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n810), .A2(new_n372), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n866), .A2(new_n733), .A3(new_n881), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n722), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1090), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n919), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1113), .A2(new_n1139), .ZN(G378));
  OAI21_X1  g0940(.A(new_n378), .B1(new_n620), .B2(new_n621), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n377), .A2(new_n642), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT55), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n378), .B(new_n1143), .C1(new_n620), .C2(new_n621), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(new_n734), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n752), .A2(new_n768), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n767), .A2(new_n409), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G68), .B2(new_n756), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n477), .B2(new_n760), .C1(new_n279), .C2(new_n770), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1152), .B(new_n1155), .C1(G107), .C2(new_n818), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n247), .A2(new_n262), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n773), .A2(G116), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1156), .A2(new_n1020), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT58), .Z(new_n1160));
  OAI221_X1 g0960(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n247), .C2(new_n262), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n785), .A2(new_n1121), .B1(G125), .B2(new_n773), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n764), .A2(new_n1118), .B1(new_n770), .B2(new_n823), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G150), .B2(new_n756), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(new_n821), .C2(new_n760), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT114), .B(KEYINPUT59), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n399), .B2(new_n767), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n736), .B1(new_n1160), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n713), .B1(new_n202), .B2(new_n810), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1151), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT116), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1150), .B1(new_n896), .B2(G330), .ZN(new_n1176));
  AND4_X1   g0976(.A1(G330), .A2(new_n899), .A3(new_n900), .A4(new_n1150), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n888), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n901), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n896), .A2(G330), .A3(new_n1150), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1175), .A3(new_n887), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1174), .B1(new_n1185), .B2(new_n919), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1112), .A2(new_n1102), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n887), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT96), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n864), .B(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1191), .A2(new_n1181), .A3(new_n885), .A4(new_n1182), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1188), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n661), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1185), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1186), .B1(new_n1195), .B2(new_n1196), .ZN(G375));
  NOR2_X1   g0997(.A1(new_n1110), .A2(new_n920), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n782), .A2(new_n1015), .B1(new_n770), .B2(new_n251), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G116), .B2(new_n759), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT117), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n247), .B(new_n1201), .C1(G97), .C2(new_n749), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n768), .B2(new_n764), .C1(new_n599), .C2(new_n752), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1203), .A2(new_n991), .A3(new_n1024), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n749), .A2(G159), .B1(G128), .B2(new_n753), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n247), .B1(new_n782), .B2(new_n821), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n770), .A2(new_n365), .B1(new_n755), .B2(new_n202), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1206), .A2(new_n1153), .A3(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(new_n823), .C2(new_n764), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n759), .B2(new_n1121), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n736), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n722), .C1(new_n734), .C2(new_n840), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n216), .B2(new_n810), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1198), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n955), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1111), .B2(new_n1216), .ZN(G381));
  NOR2_X1   g1017(.A1(G375), .A2(G378), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G381), .A2(G384), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1009), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n957), .B2(new_n981), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1223), .A2(G396), .A3(G393), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1218), .A2(new_n1219), .A3(new_n1224), .ZN(G407));
  INV_X1    g1025(.A(G213), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G343), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1218), .A2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT118), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT118), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(G213), .A3(G407), .A4(new_n1230), .ZN(G409));
  NAND2_X1  g1031(.A1(G387), .A2(G390), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(G393), .B(new_n791), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1232), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G387), .A2(KEYINPUT124), .A3(G390), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT124), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1222), .B1(new_n1221), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1233), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1186), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1187), .A2(new_n1185), .A3(new_n955), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1174), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n919), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1136), .B1(new_n1100), .B2(new_n920), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1112), .A2(new_n661), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1109), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1227), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1215), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1110), .A2(new_n1101), .A3(KEYINPUT60), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n1108), .A3(new_n661), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1214), .ZN(new_n1260));
  INV_X1    g1060(.A(G384), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT119), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1261), .A2(KEYINPUT119), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1259), .A2(KEYINPUT119), .A3(new_n1261), .A4(new_n1214), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1227), .A2(KEYINPUT122), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1227), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1269), .A3(new_n1267), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1243), .B(new_n1244), .C1(new_n1255), .C2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1255), .A2(new_n1275), .A3(new_n1266), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1255), .B2(new_n1266), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1245), .A2(new_n1254), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1227), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT121), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1273), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT121), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1255), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1266), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1227), .B(new_n1287), .C1(new_n1245), .C2(new_n1254), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT120), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  OAI211_X1 g1092(.A(KEYINPUT120), .B(new_n1292), .C1(new_n1281), .C2(new_n1287), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1286), .A2(new_n1289), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1278), .B1(new_n1294), .B2(new_n1295), .ZN(G405));
  AOI21_X1  g1096(.A(KEYINPUT127), .B1(new_n1266), .B2(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1297), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1243), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1253), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1302), .A2(KEYINPUT125), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1266), .A2(KEYINPUT127), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(KEYINPUT125), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1245), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1301), .B(new_n1306), .ZN(G402));
endmodule


