//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  AND3_X1   g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT64), .B(G238), .Z(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n222), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n203), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n249), .B1(new_n250), .B2(new_n252), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n226), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n254), .A3(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n202), .ZN(new_n262));
  INV_X1    g0062(.A(new_n258), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G1), .B2(new_n254), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(new_n202), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n259), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n277), .B(new_n278), .C1(G77), .C2(new_n273), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT67), .B(G226), .Z(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT68), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G41), .B2(G45), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n282), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n279), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT70), .B(G200), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n259), .A2(KEYINPUT9), .A3(new_n265), .A4(new_n262), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n279), .A2(new_n288), .A3(G190), .A4(new_n291), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n268), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n266), .B1(new_n292), .B2(G179), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n292), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT76), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n207), .A2(G1698), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(G226), .B2(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT73), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n278), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G238), .B1(new_n286), .B2(new_n287), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n291), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT13), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .A4(new_n291), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n307), .B1(new_n322), .B2(G169), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n301), .B(new_n306), .C1(new_n319), .C2(new_n321), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT74), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n327), .A3(new_n321), .ZN(new_n328));
  OR3_X1    g0128(.A1(new_n318), .A2(new_n327), .A3(KEYINPUT13), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n215), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n333), .B1(new_n255), .B2(new_n334), .C1(new_n252), .C2(new_n202), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n258), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(new_n258), .A3(new_n337), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n333), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n260), .A2(G1), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT12), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(KEYINPUT12), .A3(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n215), .B2(new_n264), .ZN(new_n347));
  NOR4_X1   g0147(.A1(new_n340), .A2(new_n342), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n332), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(G20), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G77), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n264), .A2(new_n334), .ZN(new_n353));
  INV_X1    g0153(.A(new_n253), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  INV_X1    g0155(.A(new_n255), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n354), .A2(new_n251), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n254), .B2(new_n334), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n352), .B(new_n353), .C1(new_n358), .C2(new_n258), .ZN(new_n359));
  OAI21_X1  g0159(.A(G244), .B1(new_n286), .B2(new_n287), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(new_n291), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n275), .A2(G232), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n273), .B(new_n362), .C1(new_n216), .C2(new_n275), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n278), .C1(G107), .C2(new_n273), .ZN(new_n364));
  AOI21_X1  g0164(.A(G169), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT71), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n352), .B1(new_n358), .B2(new_n258), .ZN(new_n367));
  INV_X1    g0167(.A(new_n353), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(new_n291), .A3(new_n360), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n301), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n361), .A2(new_n326), .A3(new_n364), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n366), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n370), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n293), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT69), .B1(new_n370), .B2(new_n376), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n377), .A2(new_n359), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n319), .B2(new_n321), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n328), .A2(new_n329), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n348), .B(new_n385), .C1(new_n386), .C2(new_n376), .ZN(new_n387));
  AND4_X1   g0187(.A1(new_n303), .A2(new_n350), .A3(new_n382), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n309), .A2(new_n310), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n389), .B2(new_n254), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n254), .A4(new_n272), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n201), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n251), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n400), .A3(new_n396), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n393), .A2(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n271), .A2(new_n254), .A3(new_n272), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n215), .B1(new_n405), .B2(new_n391), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n399), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(new_n397), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n258), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT78), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n273), .B1(G223), .B2(G1698), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n275), .A2(G226), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(new_n270), .B2(new_n208), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n290), .B1(new_n413), .B2(new_n278), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n376), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n278), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n417), .A2(new_n415), .A3(new_n291), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(G200), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n253), .A2(new_n261), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n264), .B2(new_n253), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n393), .A2(KEYINPUT77), .A3(new_n399), .A4(new_n398), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n407), .B1(new_n406), .B2(new_n397), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n258), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n410), .A2(new_n419), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n425), .B2(new_n258), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT78), .B(new_n263), .C1(new_n423), .C2(new_n424), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n431), .A2(new_n432), .A3(new_n421), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n419), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n410), .A2(new_n422), .A3(new_n427), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n414), .A2(new_n415), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n301), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n417), .A2(new_n326), .A3(new_n415), .A4(new_n291), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT79), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT79), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n414), .A2(new_n440), .A3(new_n326), .A4(new_n415), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT18), .B1(new_n435), .B2(new_n442), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n430), .B(new_n434), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n388), .A2(KEYINPUT80), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT80), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n350), .A2(new_n303), .A3(new_n382), .A4(new_n387), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n428), .B(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n433), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n435), .A2(new_n442), .A3(KEYINPUT18), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n447), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n449), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n270), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n273), .A2(G238), .A3(new_n275), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT82), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n273), .A2(new_n465), .A3(G238), .A4(new_n275), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n467), .A2(new_n282), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n282), .B(G250), .C1(G1), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(G1), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G274), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n468), .A2(new_n326), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n355), .A2(new_n351), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n263), .B(new_n351), .C1(G1), .C2(new_n270), .ZN(new_n476));
  INV_X1    g0276(.A(new_n355), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n313), .A2(new_n314), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT19), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n254), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n273), .A2(new_n254), .A3(G68), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT19), .B1(new_n356), .B2(G97), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n475), .B(new_n478), .C1(new_n487), .C2(new_n263), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n315), .B2(KEYINPUT19), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n484), .B(new_n491), .C1(new_n492), .C2(new_n479), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n474), .B1(new_n493), .B2(new_n258), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT83), .A3(new_n478), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n470), .B(new_n472), .C1(new_n467), .C2(new_n282), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n301), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n473), .A2(new_n490), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n293), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n476), .A2(new_n208), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n474), .B(new_n500), .C1(new_n493), .C2(new_n258), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n501), .C1(new_n376), .C2(new_n496), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n261), .A2(new_n217), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n476), .B2(new_n217), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n390), .B2(new_n392), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n217), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(KEYINPUT6), .A3(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n251), .A2(G77), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n505), .B1(new_n516), .B2(new_n258), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(G244), .C1(new_n310), .C2(new_n309), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  INV_X1    g0322(.A(G244), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n271), .B2(new_n272), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n522), .C1(new_n524), .C2(KEYINPUT4), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n309), .B2(new_n310), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n275), .B1(new_n526), .B2(KEYINPUT4), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n278), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT5), .B(G41), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G274), .A3(new_n471), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n278), .B1(new_n471), .B2(new_n529), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G257), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n301), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n528), .A2(new_n326), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n518), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n254), .B(G87), .C1(new_n309), .C2(new_n310), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n273), .A2(new_n540), .A3(new_n254), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT23), .A3(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT23), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n270), .A2(new_n461), .B1(new_n545), .B2(KEYINPUT85), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n254), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n254), .B2(G107), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n545), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n542), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n549), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n539), .B2(new_n541), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n544), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n258), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n209), .A2(new_n275), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n218), .A2(G1698), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n309), .C2(new_n310), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G294), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n282), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(G264), .B2(new_n532), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G190), .A3(new_n530), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n530), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n476), .A2(new_n508), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n344), .A2(G20), .A3(new_n508), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT25), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n558), .A2(new_n565), .A3(new_n567), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n534), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n528), .A2(G190), .A3(new_n533), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n517), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n573), .A2(new_n517), .A3(new_n577), .A4(new_n574), .ZN(new_n578));
  AND4_X1   g0378(.A1(new_n537), .A2(new_n572), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n522), .B(new_n254), .C1(G33), .C2(new_n217), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n263), .B1(KEYINPUT84), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n461), .A2(G20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n270), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n254), .A4(new_n522), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(KEYINPUT84), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(new_n258), .A3(new_n582), .A4(new_n585), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n476), .A2(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n351), .A2(new_n461), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n532), .A2(G270), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n275), .A2(G257), .ZN(new_n597));
  INV_X1    g0397(.A(G264), .ZN(new_n598));
  OAI221_X1 g0398(.A(new_n597), .B1(new_n598), .B2(new_n275), .C1(new_n309), .C2(new_n310), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n389), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n601), .A3(new_n278), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n596), .A2(new_n530), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n595), .A2(KEYINPUT21), .A3(G169), .A4(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n586), .A2(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n376), .C2(new_n603), .ZN(new_n607));
  INV_X1    g0407(.A(new_n603), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n595), .A2(G179), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(G169), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n604), .A2(new_n607), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(G169), .B1(new_n564), .B2(new_n530), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n598), .B(new_n278), .C1(new_n471), .C2(new_n529), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n615), .A2(new_n563), .A3(G179), .A4(new_n531), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n263), .B1(new_n552), .B2(new_n556), .ZN(new_n618));
  INV_X1    g0418(.A(new_n571), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT86), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT86), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n617), .B(new_n622), .C1(new_n618), .C2(new_n619), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n613), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n459), .A2(new_n503), .A3(new_n579), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n537), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n498), .A2(new_n626), .A3(new_n502), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n497), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n301), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(new_n473), .A3(new_n488), .A4(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n502), .A4(new_n626), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n632), .A2(new_n502), .A3(new_n572), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n576), .A2(new_n537), .A3(new_n578), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n604), .A2(new_n612), .A3(new_n609), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT88), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n604), .A2(new_n609), .A3(new_n612), .A4(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n620), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n638), .B(new_n640), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n636), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n459), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n375), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n349), .A2(new_n332), .B1(new_n387), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n434), .A2(new_n430), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n456), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n299), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n302), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n649), .A2(new_n655), .ZN(G369));
  NOR2_X1   g0456(.A1(new_n260), .A2(G20), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n284), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  INV_X1    g0460(.A(G213), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n645), .A2(new_n605), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n641), .ZN(new_n665));
  INV_X1    g0465(.A(new_n663), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n665), .A2(new_n607), .B1(new_n595), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n621), .A2(new_n623), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n666), .B1(new_n618), .B2(new_n619), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n572), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n620), .B2(new_n663), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n641), .A2(new_n663), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n620), .B2(new_n666), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n678), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n223), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G1), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n479), .A2(new_n461), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n230), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n666), .B1(new_n636), .B2(new_n647), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT91), .B1(new_n690), .B2(KEYINPUT29), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n646), .B1(new_n642), .B2(new_n644), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n692), .A2(new_n639), .A3(new_n637), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n663), .B1(new_n693), .B2(new_n635), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n639), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n576), .A2(KEYINPUT92), .A3(new_n537), .A4(new_n578), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n673), .A2(new_n665), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n638), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n632), .A2(new_n502), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n626), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n503), .A2(new_n633), .A3(new_n626), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n703), .A2(new_n706), .A3(new_n632), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n691), .A2(new_n697), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n496), .A2(new_n534), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n603), .A2(new_n326), .A3(new_n563), .A4(new_n615), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n608), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n496), .A3(new_n534), .A4(new_n566), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT90), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n712), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT90), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n721), .A3(new_n717), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n715), .A2(new_n717), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n663), .B1(new_n726), .B2(new_n720), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n579), .A2(new_n624), .A3(new_n503), .A4(new_n663), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(KEYINPUT31), .ZN(new_n729));
  OAI21_X1  g0529(.A(G330), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n689), .B1(new_n731), .B2(G1), .ZN(G364));
  XNOR2_X1  g0532(.A(new_n668), .B(KEYINPUT89), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n670), .A2(new_n671), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n686), .B1(G45), .B2(new_n657), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n683), .A2(new_n273), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n229), .A2(new_n469), .A3(G50), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(new_n247), .C2(new_n469), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n683), .A2(new_n389), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G355), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n741), .B(new_n743), .C1(G116), .C2(new_n223), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n226), .B1(G20), .B2(new_n301), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n737), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n254), .A2(new_n326), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n383), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G326), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n326), .A2(new_n383), .A3(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n753), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G322), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G311), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n254), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n293), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n376), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G303), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n763), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n752), .A2(new_n376), .A3(G200), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  OAI221_X1 g0574(.A(new_n389), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n768), .A2(G190), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(G283), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n762), .A2(new_n766), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n759), .A2(new_n217), .B1(new_n334), .B2(new_n764), .ZN(new_n779));
  INV_X1    g0579(.A(new_n776), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n508), .ZN(new_n781));
  INV_X1    g0581(.A(new_n773), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n779), .B(new_n781), .C1(G68), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n389), .B1(new_n769), .B2(G87), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n786));
  INV_X1    g0586(.A(new_n754), .ZN(new_n787));
  INV_X1    g0587(.A(new_n771), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n202), .B1(new_n789), .B2(KEYINPUT32), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(KEYINPUT32), .B2(new_n789), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n761), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n206), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n778), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  INV_X1    g0596(.A(new_n747), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n750), .B1(new_n751), .B2(new_n796), .C1(new_n733), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n738), .A2(new_n798), .ZN(G396));
  NOR2_X1   g0599(.A1(new_n359), .A2(new_n663), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n375), .A2(new_n380), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n366), .A2(new_n373), .A3(new_n800), .A4(new_n374), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n694), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(new_n730), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n737), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n761), .B1(new_n782), .B2(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n787), .C1(new_n810), .C2(new_n764), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT34), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n776), .A2(G68), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n206), .B2(new_n759), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  INV_X1    g0617(.A(new_n769), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n273), .B1(new_n817), .B2(new_n771), .C1(new_n818), .C2(new_n202), .ZN(new_n819));
  OR4_X1    g0619(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n773), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n759), .A2(new_n217), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n787), .A2(new_n600), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(G294), .C2(new_n761), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n389), .B1(new_n771), .B2(new_n826), .C1(new_n461), .C2(new_n764), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G107), .B2(new_n769), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n828), .C1(new_n208), .C2(new_n780), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n820), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n751), .A2(new_n746), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n830), .A2(new_n748), .B1(new_n334), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n736), .C1(new_n746), .C2(new_n804), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n807), .A2(new_n834), .ZN(G384));
  NAND2_X1  g0635(.A1(new_n435), .A2(new_n442), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n435), .A2(new_n662), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n428), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n399), .B1(new_n406), .B2(new_n397), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n258), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n422), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n442), .B2(new_n662), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n844), .A2(new_n428), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n839), .B1(new_n845), .B2(new_n838), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT96), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n843), .A2(new_n662), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(new_n451), .C2(new_n456), .ZN(new_n849));
  INV_X1    g0649(.A(new_n848), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT96), .B1(new_n445), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT38), .B(new_n846), .C1(new_n849), .C2(new_n851), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n836), .A2(new_n837), .A3(new_n428), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(new_n838), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n837), .B1(new_n451), .B2(new_n456), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n350), .A2(new_n666), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n856), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n376), .B1(new_n328), .B2(new_n329), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n866), .A2(new_n349), .A3(new_n384), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n349), .B(new_n666), .C1(new_n332), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n349), .A2(new_n666), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n330), .A2(new_n323), .A3(new_n324), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n387), .B(new_n869), .C1(new_n870), .C2(new_n348), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n650), .A2(new_n663), .ZN(new_n873));
  INV_X1    g0673(.A(new_n804), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n694), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n851), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n445), .A2(KEYINPUT96), .A3(new_n850), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n878), .B2(new_n846), .ZN(new_n879));
  INV_X1    g0679(.A(new_n855), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n872), .B(new_n875), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n456), .A2(new_n662), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n865), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n459), .A2(new_n691), .A3(new_n709), .A4(new_n697), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n655), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n883), .B(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n855), .A2(new_n860), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n874), .B1(new_n868), .B2(new_n871), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n729), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT98), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n888), .B(KEYINPUT98), .C1(new_n729), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT40), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT97), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT40), .B1(new_n890), .B2(new_n896), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(new_n879), .C2(new_n880), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n729), .A2(new_n889), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n459), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n900), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n886), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n284), .B2(new_n657), .ZN(new_n907));
  OAI211_X1 g0707(.A(G20), .B(new_n227), .C1(new_n513), .C2(KEYINPUT35), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n461), .B(new_n908), .C1(KEYINPUT35), .C2(new_n513), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT36), .Z(new_n910));
  OAI21_X1  g0710(.A(G77), .B1(new_n206), .B2(new_n215), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n230), .A2(new_n911), .B1(G50), .B2(new_n215), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n260), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n907), .A2(new_n910), .A3(new_n913), .ZN(G367));
  OAI21_X1  g0714(.A(new_n704), .B1(new_n501), .B2(new_n663), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n632), .A2(new_n501), .A3(new_n663), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT43), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n517), .A2(new_n663), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n920), .B(new_n673), .C1(new_n699), .C2(new_n700), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT99), .B1(new_n921), .B2(new_n626), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT99), .ZN(new_n923));
  INV_X1    g0723(.A(new_n920), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n701), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n537), .C1(new_n925), .C2(new_n673), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n926), .A3(new_n663), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n675), .A2(new_n679), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT42), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n920), .B1(new_n699), .B2(new_n700), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n927), .A2(KEYINPUT100), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT100), .B1(new_n927), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n919), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT101), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n915), .A2(new_n918), .A3(new_n916), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT101), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n919), .C1(new_n934), .C2(new_n935), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT102), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n930), .B1(new_n626), .B2(new_n666), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n677), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n942), .A2(new_n943), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(KEYINPUT103), .A3(new_n946), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n950), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT103), .B1(new_n944), .B2(new_n946), .ZN(new_n954));
  INV_X1    g0754(.A(new_n946), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n948), .B(new_n955), .C1(new_n942), .C2(new_n943), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n681), .A2(new_n945), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n681), .A2(new_n945), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n960));
  OR2_X1    g0760(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n678), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n677), .A2(new_n959), .A3(new_n962), .A4(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n679), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n680), .B(KEYINPUT105), .C1(new_n676), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(KEYINPUT105), .B2(new_n680), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n734), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n731), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n731), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n684), .B(KEYINPUT41), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n657), .A2(G45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(G1), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n952), .A2(new_n957), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n389), .B1(new_n771), .B2(new_n982), .C1(new_n821), .C2(new_n764), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n761), .A2(G303), .B1(G107), .B2(new_n758), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n826), .B2(new_n787), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G97), .C2(new_n776), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n769), .A2(G116), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(new_n756), .C2(new_n773), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT107), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n764), .A2(new_n202), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n759), .A2(new_n215), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n793), .A2(new_n250), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G143), .C2(new_n754), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n273), .B1(new_n771), .B2(new_n809), .C1(new_n773), .C2(new_n810), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G58), .B2(new_n769), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n334), .C2(new_n780), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n737), .B1(new_n999), .B2(new_n748), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n739), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n749), .B1(new_n223), .B2(new_n477), .C1(new_n240), .C2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(new_n797), .C2(new_n917), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n981), .A2(new_n1003), .ZN(G387));
  OR2_X1    g0804(.A1(new_n971), .A2(new_n731), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n684), .A3(new_n972), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n971), .A2(new_n978), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1001), .B1(new_n237), .B2(G45), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n687), .B2(new_n742), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n354), .A2(new_n202), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n687), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1011), .B(new_n469), .C1(KEYINPUT50), .C2(new_n1010), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G68), .B2(G77), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n223), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n737), .B1(new_n1014), .B2(new_n749), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n761), .B1(new_n782), .B2(G311), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n754), .A2(G322), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n600), .C2(new_n764), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n821), .B2(new_n759), .C1(new_n756), .C2(new_n818), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n788), .A2(G326), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n273), .B1(new_n776), .B2(G116), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n202), .A2(new_n793), .B1(new_n787), .B2(new_n810), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n477), .A2(new_n759), .B1(new_n253), .B2(new_n773), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n389), .B1(new_n788), .B2(G150), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n818), .B2(new_n334), .C1(new_n217), .C2(new_n780), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT109), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1028), .B(new_n1029), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .C1(new_n215), .C2(new_n764), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1016), .B1(new_n676), .B2(new_n797), .C1(new_n1035), .C2(new_n751), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1006), .A2(new_n1007), .A3(new_n1036), .ZN(G393));
  INV_X1    g0837(.A(KEYINPUT110), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n966), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n972), .C1(new_n967), .C2(KEYINPUT110), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n967), .A2(new_n972), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n684), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n945), .A2(new_n747), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n223), .A2(new_n217), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n749), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n244), .C2(new_n739), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n389), .B1(new_n764), .B2(new_n756), .C1(new_n759), .C2(new_n461), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1047), .B(new_n781), .C1(G303), .C2(new_n782), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n769), .A2(G283), .B1(G322), .B2(new_n788), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  AOI22_X1  g0850(.A1(G311), .A2(new_n761), .B1(new_n754), .B2(G317), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1052));
  XNOR2_X1  g0852(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT115), .Z(new_n1055));
  AOI22_X1  g0855(.A1(G150), .A2(new_n754), .B1(new_n761), .B2(G159), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G68), .A2(new_n769), .B1(new_n776), .B2(G87), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n773), .A2(new_n202), .B1(new_n764), .B2(new_n253), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT112), .Z(new_n1061));
  NOR2_X1   g0861(.A1(new_n759), .A2(new_n334), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n389), .B(new_n1062), .C1(G143), .C2(new_n788), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n751), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1043), .A2(new_n737), .A3(new_n1046), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1039), .B1(new_n967), .B2(KEYINPUT110), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n978), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1042), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G390));
  NAND3_X1  g0870(.A1(new_n459), .A2(G330), .A3(new_n902), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n884), .A2(new_n655), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n804), .A2(G330), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n872), .B(new_n1074), .C1(new_n729), .C2(new_n889), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n727), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1073), .B1(new_n1078), .B2(new_n724), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1075), .B1(new_n1079), .B2(new_n872), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n875), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n872), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n868), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n901), .B2(new_n1073), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n708), .A2(new_n663), .A3(new_n804), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n872), .B(new_n1074), .C1(new_n725), .C2(new_n729), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n873), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1072), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1075), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n864), .B1(new_n875), .B2(new_n872), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT39), .B1(new_n855), .B2(new_n860), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1085), .B1(new_n1087), .B2(new_n873), .ZN(new_n1099));
  OR3_X1    g0899(.A1(new_n887), .A2(new_n1099), .A3(new_n864), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1093), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1094), .B1(new_n856), .B2(new_n863), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n887), .A2(new_n1099), .A3(new_n864), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1088), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1088), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1098), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1075), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n1092), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n684), .C1(new_n1110), .C2(new_n1092), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n978), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n745), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n737), .B1(new_n832), .B2(new_n253), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT118), .ZN(new_n1118));
  INV_X1    g0918(.A(G128), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1119), .A2(new_n787), .B1(new_n793), .B2(new_n817), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT54), .B(G143), .Z(new_n1121));
  AOI21_X1  g0921(.A(new_n389), .B1(new_n765), .B2(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n809), .B2(new_n773), .C1(new_n780), .C2(new_n202), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1120), .B(new_n1123), .C1(G159), .C2(new_n758), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n769), .A2(G150), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT53), .Z(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1124), .B(new_n1126), .C1(new_n1127), .C2(new_n771), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n787), .A2(new_n821), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1062), .B(new_n1129), .C1(G116), .C2(new_n761), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n769), .A2(G87), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n389), .B1(new_n771), .B2(new_n756), .C1(new_n773), .C2(new_n508), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G97), .B2(new_n765), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .A4(new_n815), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1118), .B1(new_n1135), .B2(new_n748), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT119), .Z(new_n1137));
  NAND2_X1  g0937(.A1(new_n1116), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1114), .A2(new_n1115), .A3(new_n1138), .ZN(G378));
  NAND2_X1  g0939(.A1(new_n900), .A2(G330), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n883), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n303), .B(KEYINPUT55), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n266), .A2(new_n662), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT56), .Z(new_n1144));
  XOR2_X1   g0944(.A(new_n1142), .B(new_n1144), .Z(new_n1145));
  AOI21_X1  g0945(.A(new_n671), .B1(new_n895), .B2(new_n899), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n865), .A2(new_n881), .A3(new_n882), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1141), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1145), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1148), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1113), .A2(new_n1072), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n685), .B1(new_n1154), .B2(KEYINPUT57), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n884), .A2(new_n655), .A3(new_n1071), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1141), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1145), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1156), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1111), .B1(new_n1110), .B2(new_n1092), .ZN(new_n1164));
  AOI211_X1 g0964(.A(KEYINPUT117), .B(new_n1091), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1072), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1153), .A2(new_n1149), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT122), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n1156), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1155), .A2(new_n1163), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1145), .A2(new_n745), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n389), .B1(new_n821), .B2(new_n771), .C1(new_n780), .C2(new_n206), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G41), .B(new_n1173), .C1(G77), .C2(new_n769), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT120), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n508), .A2(new_n793), .B1(new_n787), .B2(new_n461), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n992), .B(new_n1176), .C1(G97), .C2(new_n782), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n477), .C2(new_n764), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n759), .A2(new_n250), .B1(new_n773), .B2(new_n817), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1127), .A2(new_n787), .B1(new_n793), .B2(new_n1119), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n769), .C2(new_n1121), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n809), .B2(new_n764), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT59), .Z(new_n1185));
  AOI21_X1  g0985(.A(G41), .B1(new_n776), .B2(G159), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT121), .B(G124), .Z(new_n1187));
  AOI21_X1  g0987(.A(G33), .B1(new_n788), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n202), .B1(new_n309), .B2(G41), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1180), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n748), .B1(new_n202), .B2(new_n832), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1172), .A2(new_n736), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1167), .B2(new_n978), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(new_n1196), .ZN(G375));
  AND2_X1   g0997(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1157), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n974), .A3(new_n1091), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1085), .A2(new_n745), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n793), .A2(new_n809), .B1(new_n202), .B2(new_n759), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G132), .B2(new_n754), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n782), .A2(new_n1121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n769), .A2(G159), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n273), .B1(new_n771), .B2(new_n1119), .C1(new_n250), .C2(new_n764), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G58), .B2(new_n776), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n761), .A2(G283), .B1(new_n355), .B2(new_n758), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n756), .B2(new_n787), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n389), .B1(new_n764), .B2(new_n508), .C1(new_n461), .C2(new_n773), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G77), .B2(new_n776), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n217), .C2(new_n818), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n771), .A2(new_n600), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1208), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1216), .A2(new_n748), .B1(new_n215), .B2(new_n832), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1201), .A2(new_n736), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1090), .B2(new_n978), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(G381));
  NAND3_X1  g1020(.A1(new_n981), .A2(new_n1003), .A3(new_n1069), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1221), .A2(G396), .A3(G393), .ZN(new_n1222));
  INV_X1    g1022(.A(G384), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1219), .A4(new_n1200), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT123), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1114), .A2(new_n1196), .A3(new_n1115), .A4(new_n1138), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1169), .B1(new_n1168), .B2(new_n1156), .ZN(new_n1227));
  AOI211_X1 g1027(.A(KEYINPUT122), .B(KEYINPUT57), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1226), .B1(new_n1229), .B2(new_n1155), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(KEYINPUT123), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(new_n1230), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  NOR2_X1   g1034(.A1(new_n661), .A2(G343), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1226), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1154), .A2(new_n974), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n684), .B(new_n1091), .C1(new_n1199), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT60), .B1(new_n1198), .B2(new_n1157), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1219), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(new_n1223), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1223), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1196), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1229), .B2(new_n1155), .ZN(new_n1248));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1238), .B(new_n1246), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  AND4_X1   g1053(.A1(new_n1253), .A2(new_n1245), .A3(G2897), .A4(new_n1235), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1245), .A2(new_n1253), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G2897), .B(new_n1235), .C1(new_n1245), .C2(new_n1253), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1249), .B1(new_n1171), .B2(new_n1196), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1237), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1259), .A2(new_n1226), .B1(new_n661), .B2(G343), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1238), .A4(new_n1246), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1251), .A2(new_n1252), .A3(new_n1261), .A4(new_n1264), .ZN(new_n1265));
  XOR2_X1   g1065(.A(G393), .B(G396), .Z(new_n1266));
  NAND2_X1  g1066(.A1(new_n1221), .A2(KEYINPUT126), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1069), .B1(new_n981), .B2(new_n1003), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1266), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(KEYINPUT126), .A3(new_n1221), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1261), .A2(new_n1276), .A3(new_n1252), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT124), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1258), .A2(new_n1260), .A3(new_n1245), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(KEYINPUT63), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1250), .A2(KEYINPUT124), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1277), .A2(new_n1280), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1275), .A2(new_n1284), .ZN(G405));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1273), .B(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1258), .A2(new_n1230), .A3(new_n1246), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1245), .B1(new_n1233), .B2(new_n1262), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1288), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1274), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(G402));
endmodule


