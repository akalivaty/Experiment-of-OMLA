//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT36), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT36), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT32), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G134gat), .ZN(new_n213));
  INV_X1    g012(.A(G134gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G127gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT68), .B1(new_n214), .B2(G127gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n211), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n213), .A2(new_n215), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n232));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n240), .A2(new_n226), .A3(KEYINPUT64), .A4(new_n227), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n230), .A2(new_n236), .A3(new_n237), .A4(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n243));
  INV_X1    g042(.A(new_n227), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n244), .B1(new_n247), .B2(new_n224), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n238), .A2(new_n249), .A3(new_n239), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n238), .B2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n243), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n242), .B1(new_n253), .B2(new_n237), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n231), .A2(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n238), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(new_n231), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT67), .B1(new_n224), .B2(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n247), .B(new_n261), .C1(new_n262), .C2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n262), .A3(KEYINPUT28), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n222), .B1(new_n254), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n259), .ZN(new_n272));
  INV_X1    g071(.A(new_n246), .ZN(new_n273));
  NAND2_X1  g072(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n261), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(G183gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT28), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n266), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n272), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n224), .A3(new_n274), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n229), .A2(new_n249), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n227), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n236), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT25), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n220), .A2(new_n211), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n214), .A2(G127gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n212), .A2(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n217), .B1(new_n293), .B2(KEYINPUT68), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n294), .B2(new_n211), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n283), .A2(new_n289), .A3(new_n295), .A4(new_n242), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n271), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT69), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n268), .A2(new_n296), .A3(new_n299), .A4(new_n271), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n206), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT33), .B1(new_n298), .B2(new_n300), .ZN(new_n302));
  XOR2_X1   g101(.A(G15gat), .B(G43gat), .Z(new_n303));
  XNOR2_X1  g102(.A(G71gat), .B(G99gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  AOI221_X4 g106(.A(new_n206), .B1(KEYINPUT33), .B2(new_n305), .C1(new_n298), .C2(new_n300), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n268), .A2(new_n296), .ZN(new_n311));
  INV_X1    g110(.A(new_n271), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g112(.A(new_n271), .B(new_n309), .C1(new_n268), .C2(new_n296), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n307), .A2(new_n308), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n300), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT33), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n301), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n308), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n315), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n204), .B(new_n205), .C1(new_n317), .C2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n316), .B1(new_n307), .B2(new_n308), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n323), .A3(new_n315), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT36), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT71), .A4(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n332), .A2(new_n334), .B1(KEYINPUT2), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n335), .ZN(new_n337));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT74), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G155gat), .B(G162gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT74), .B(new_n344), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n295), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT39), .B1(new_n352), .B2(KEYINPUT84), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(KEYINPUT84), .B2(new_n352), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n343), .A2(KEYINPUT3), .A3(new_n348), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n295), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n343), .A2(new_n348), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n359), .A2(new_n295), .A3(KEYINPUT4), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n222), .B2(new_n349), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(new_n351), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n222), .A2(new_n361), .A3(new_n349), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT4), .B1(new_n359), .B2(new_n295), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n357), .A2(new_n295), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n356), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT82), .B1(new_n370), .B2(new_n351), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT39), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n370), .A2(KEYINPUT82), .A3(new_n351), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(KEYINPUT81), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT83), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT39), .B1(new_n371), .B2(new_n366), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(new_n382), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n372), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  AND2_X1   g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n254), .B2(new_n267), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n399), .A2(new_n400), .B1(G211gat), .B2(G218gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n405), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n283), .A2(new_n289), .A3(new_n242), .A4(new_n395), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n398), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n398), .B2(new_n410), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT73), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(KEYINPUT73), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n393), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n410), .ZN(new_n417));
  INV_X1    g216(.A(new_n409), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT73), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n409), .A3(new_n410), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n393), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n393), .C1(new_n413), .C2(new_n415), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n365), .B1(new_n369), .B2(new_n356), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n222), .A2(KEYINPUT75), .A3(new_n361), .A4(new_n349), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n368), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n359), .B(new_n295), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n365), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT5), .B1(new_n368), .B2(new_n367), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n382), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n425), .A2(new_n427), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT40), .B(new_n372), .C1(new_n384), .C2(new_n387), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n390), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n356), .A2(new_n396), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n418), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT29), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n407), .A2(KEYINPUT79), .A3(new_n408), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT3), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(new_n349), .ZN(new_n450));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n355), .B1(new_n418), .B2(KEYINPUT29), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n359), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n444), .B2(new_n418), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G22gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(KEYINPUT80), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT80), .B1(new_n455), .B2(new_n456), .ZN(new_n465));
  INV_X1    g264(.A(new_n462), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n464), .A2(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n432), .A2(new_n435), .B1(new_n428), .B2(new_n437), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n381), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT78), .B1(new_n470), .B2(KEYINPUT6), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NOR4_X1   g272(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n381), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n413), .B2(new_n415), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n422), .A2(KEYINPUT37), .A3(new_n414), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n423), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT38), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT6), .B1(new_n469), .B2(new_n381), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n440), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n423), .B1(new_n422), .B2(new_n414), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n476), .B1(new_n419), .B2(new_n421), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n484), .A2(KEYINPUT38), .A3(new_n393), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n485), .B2(new_n477), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n475), .A2(new_n480), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n443), .A2(new_n468), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n425), .A2(new_n427), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT77), .ZN(new_n490));
  INV_X1    g289(.A(new_n381), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n490), .B(new_n473), .C1(new_n439), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n439), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n481), .A2(new_n490), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n474), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n472), .B1(new_n493), .B2(new_n473), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n489), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n468), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n330), .A2(new_n488), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n468), .A2(new_n327), .A3(new_n326), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT35), .B1(new_n475), .B2(new_n482), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n317), .A2(new_n324), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n489), .A4(new_n468), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G134gat), .B(G162gat), .Z(new_n511));
  AND2_X1   g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT41), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n511), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT95), .ZN(new_n515));
  NOR2_X1   g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  XOR2_X1   g317(.A(G43gat), .B(G50gat), .Z(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT86), .B(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT87), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n522), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n518), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n520), .A2(new_n528), .A3(new_n523), .A4(new_n524), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  INV_X1    g335(.A(G85gat), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(KEYINPUT8), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G99gat), .B(G106gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(new_n533), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n540), .A2(new_n541), .ZN(new_n545));
  INV_X1    g344(.A(new_n541), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n535), .B2(new_n539), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n530), .A2(new_n548), .B1(KEYINPUT41), .B2(new_n512), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n544), .B1(new_n543), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g350(.A(G190gat), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n543), .A2(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n225), .ZN(new_n556));
  INV_X1    g355(.A(G218gat), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n515), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G218gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n514), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G64gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n576));
  AND2_X1   g375(.A1(G57gat), .A2(G64gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n571), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G127gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT16), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n585), .B1(new_n589), .B2(KEYINPUT89), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n584), .A2(G1gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n596));
  AOI21_X1  g395(.A(G8gat), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n575), .A2(new_n578), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT93), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n575), .A2(new_n605), .A3(new_n578), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n583), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n609), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n567), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n541), .A2(KEYINPUT96), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n548), .A2(new_n579), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n575), .A2(new_n578), .A3(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n542), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n604), .A2(new_n548), .A3(KEYINPUT10), .A4(new_n606), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n621), .B2(new_n622), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n617), .B2(new_n619), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n630), .A4(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n635), .B1(new_n629), .B2(new_n631), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n615), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n532), .A2(new_n602), .A3(new_n533), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n530), .A2(new_n601), .A3(new_n598), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n646), .A2(KEYINPUT18), .A3(new_n647), .A4(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n602), .A2(new_n527), .A3(new_n529), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n647), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n648), .B(KEYINPUT13), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT91), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G113gat), .B(G141gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G169gat), .B(G197gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT12), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n660), .B(new_n666), .C1(new_n651), .C2(new_n657), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n615), .B2(new_n643), .ZN(new_n672));
  AND4_X1   g471(.A1(new_n510), .A2(new_n645), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n496), .A2(new_n499), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  INV_X1    g475(.A(new_n489), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n673), .A2(new_n686), .A3(new_n507), .ZN(new_n687));
  INV_X1    g486(.A(new_n330), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n501), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NOR3_X1   g492(.A1(new_n558), .A2(new_n559), .A3(new_n566), .ZN(new_n694));
  INV_X1    g493(.A(new_n515), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n562), .B2(new_n563), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n670), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n614), .A2(new_n698), .A3(new_n643), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n510), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n674), .A3(new_n521), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n510), .B2(new_n697), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n697), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n502), .A2(KEYINPUT103), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n500), .A2(new_n501), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n706), .A2(new_n330), .A3(new_n488), .A4(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n709), .B2(new_n509), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n699), .B(KEYINPUT102), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n674), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n702), .B1(new_n715), .B2(new_n521), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n522), .A3(new_n677), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT105), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT104), .Z(new_n721));
  AOI21_X1  g520(.A(new_n522), .B1(new_n713), .B2(new_n677), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(G1329gat));
  NAND2_X1  g522(.A1(new_n713), .A2(new_n688), .ZN(new_n724));
  INV_X1    g523(.A(new_n507), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(G43gat), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n724), .A2(G43gat), .B1(new_n700), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n501), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT48), .B1(new_n730), .B2(KEYINPUT106), .ZN(new_n731));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n700), .A2(new_n732), .A3(new_n501), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n731), .B(new_n734), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n709), .A2(new_n509), .ZN(new_n736));
  INV_X1    g535(.A(new_n643), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n615), .A2(new_n670), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n674), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT107), .B(G57gat), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n677), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT49), .B(G64gat), .Z(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n739), .A2(new_n747), .A3(new_n507), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n739), .A2(new_n688), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n747), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n739), .A2(new_n501), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(G78gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1335gat));
  INV_X1    g554(.A(new_n614), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n698), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n737), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n704), .B2(new_n710), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(new_n758), .C1(new_n704), .C2(new_n710), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n674), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n757), .A2(new_n567), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n736), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n643), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n674), .A2(new_n537), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n759), .B2(new_n489), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n489), .A2(G92gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n643), .B(new_n774), .C1(new_n767), .C2(new_n768), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n677), .A3(new_n762), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n775), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n779), .B2(KEYINPUT52), .ZN(new_n780));
  INV_X1    g579(.A(new_n775), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n777), .B2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n782), .A2(new_n783), .A3(new_n773), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n776), .B1(new_n780), .B2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n763), .B2(new_n330), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n725), .A2(G99gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n769), .B2(new_n787), .ZN(G1338gat));
  OR2_X1    g587(.A1(new_n468), .A2(G106gat), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n769), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(G106gat), .B1(new_n759), .B2(new_n468), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n790), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n760), .A2(new_n501), .A3(new_n762), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(G106gat), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n796), .B2(new_n791), .ZN(G1339gat));
  OAI21_X1  g596(.A(new_n635), .B1(new_n625), .B2(KEYINPUT54), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n626), .B(new_n628), .C1(new_n621), .C2(new_n622), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n623), .B2(new_n624), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n621), .A2(KEYINPUT112), .A3(new_n628), .A4(new_n622), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n798), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(KEYINPUT55), .B1(new_n639), .B2(new_n640), .ZN(new_n808));
  INV_X1    g607(.A(new_n666), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n646), .A2(new_n647), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n810), .A2(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n658), .A2(new_n809), .B1(new_n665), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n806), .A2(KEYINPUT54), .A3(new_n627), .A4(new_n630), .ZN(new_n813));
  INV_X1    g612(.A(new_n798), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n697), .A2(new_n808), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n670), .A2(new_n808), .A3(new_n817), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n643), .A2(new_n812), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n567), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n614), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n615), .A2(new_n670), .A3(new_n643), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n764), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n504), .A2(new_n677), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n670), .ZN(new_n831));
  INV_X1    g630(.A(new_n826), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n833), .A3(new_n468), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n826), .B2(new_n501), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n764), .A2(new_n725), .A3(new_n677), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n698), .A2(new_n209), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(G1340gat));
  AOI21_X1  g640(.A(G120gat), .B1(new_n830), .B2(new_n643), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n737), .A2(new_n207), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n839), .B2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n838), .B2(new_n756), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n212), .A3(new_n614), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  NOR3_X1   g646(.A1(new_n829), .A2(G134gat), .A3(new_n567), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n838), .B2(new_n567), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1343gat));
  NAND2_X1  g650(.A1(new_n330), .A2(new_n501), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n827), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n827), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n698), .A2(G141gat), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n855), .A2(new_n857), .A3(new_n489), .A4(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n677), .B1(new_n854), .B2(KEYINPUT119), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n858), .A4(new_n857), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n688), .A2(new_n764), .A3(new_n677), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n468), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n670), .A2(new_n808), .ZN(new_n870));
  AOI211_X1 g669(.A(KEYINPUT114), .B(new_n798), .C1(new_n802), .C2(new_n806), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n813), .B2(new_n814), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n874));
  NOR3_X1   g673(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n821), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n821), .B(KEYINPUT116), .C1(new_n870), .C2(new_n875), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n567), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n614), .B1(new_n880), .B2(new_n819), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n867), .B(new_n869), .C1(new_n881), .C2(new_n825), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n868), .B1(new_n826), .B2(new_n468), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n825), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n697), .B1(new_n876), .B2(new_n877), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n818), .A2(new_n808), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n886), .A2(new_n879), .B1(new_n697), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n888), .B2(new_n614), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n867), .B1(new_n889), .B2(new_n869), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n670), .B(new_n866), .C1(new_n884), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  NOR4_X1   g691(.A1(new_n854), .A2(G141gat), .A3(new_n677), .A4(new_n698), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n891), .B2(G141gat), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n865), .A2(new_n892), .B1(new_n862), .B2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n866), .B1(new_n884), .B2(new_n890), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(G148gat), .C1(new_n897), .C2(new_n737), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n645), .A2(new_n698), .A3(new_n672), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n868), .B(new_n501), .C1(new_n899), .C2(new_n881), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n826), .B2(new_n468), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n866), .A2(new_n643), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n333), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n898), .B1(new_n904), .B2(new_n896), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n863), .A2(new_n333), .A3(new_n643), .A4(new_n857), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1345gat));
  OAI211_X1 g706(.A(new_n614), .B(new_n866), .C1(new_n884), .C2(new_n890), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G155gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n756), .A2(G155gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n863), .A2(new_n857), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT121), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n909), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n897), .B2(new_n567), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n567), .A2(G162gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n863), .A2(new_n857), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n826), .A2(new_n674), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(new_n677), .A3(new_n468), .A4(new_n507), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(G169gat), .A3(new_n698), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT122), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n674), .A2(new_n489), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n725), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n836), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n698), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(G1348gat));
  OAI21_X1  g729(.A(G176gat), .B1(new_n928), .B2(new_n737), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n737), .A2(G176gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n922), .B2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n928), .B2(new_n756), .ZN(new_n934));
  NAND2_X1  g733(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n614), .A2(new_n262), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n922), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1350gat));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n725), .B(new_n926), .C1(new_n834), .C2(new_n835), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n697), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT61), .B(new_n225), .C1(new_n947), .C2(new_n697), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n697), .A2(new_n247), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n922), .B2(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n688), .A2(new_n926), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n902), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n698), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n852), .A2(new_n489), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n921), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n921), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n670), .A3(new_n961), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n954), .A2(new_n956), .B1(new_n955), .B2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n954), .A2(new_n643), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n958), .A2(G204gat), .A3(new_n737), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  NAND4_X1  g767(.A1(new_n900), .A2(new_n614), .A3(new_n901), .A4(new_n953), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n959), .A2(new_n961), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n756), .A2(G211gat), .ZN(new_n973));
  OAI22_X1  g772(.A1(new_n970), .A2(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n697), .A3(new_n961), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n557), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n978), .A3(new_n557), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n697), .A2(G218gat), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  AOI22_X1  g780(.A1(new_n977), .A2(new_n979), .B1(new_n954), .B2(new_n981), .ZN(G1355gat));
endmodule


