

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n661, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771;

  INV_X1 U365 ( .A(n661), .ZN(n348) );
  INV_X1 U366 ( .A(KEYINPUT56), .ZN(n346) );
  INV_X1 U367 ( .A(n737), .ZN(n350) );
  INV_X1 U368 ( .A(n737), .ZN(n353) );
  INV_X1 U369 ( .A(n658), .ZN(n352) );
  XNOR2_X1 U370 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U371 ( .A(n646), .B(KEYINPUT119), .ZN(n647) );
  XOR2_X1 U372 ( .A(n657), .B(KEYINPUT62), .Z(n658) );
  INV_X1 U373 ( .A(KEYINPUT33), .ZN(n356) );
  NAND2_X1 U374 ( .A1(n540), .A2(G214), .ZN(n703) );
  BUF_X1 U375 ( .A(n530), .Z(n380) );
  XNOR2_X1 U376 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n446) );
  INV_X1 U377 ( .A(KEYINPUT65), .ZN(n484) );
  XNOR2_X2 U378 ( .A(n591), .B(n366), .ZN(n369) );
  XNOR2_X2 U379 ( .A(n465), .B(n464), .ZN(n752) );
  NOR2_X2 U380 ( .A1(G902), .A2(n733), .ZN(n474) );
  NOR2_X2 U381 ( .A1(n615), .A2(n405), .ZN(n616) );
  AND2_X2 U382 ( .A1(n628), .A2(n627), .ZN(n755) );
  XNOR2_X2 U383 ( .A(n409), .B(n609), .ZN(n716) );
  AND2_X2 U384 ( .A1(n587), .A2(n688), .ZN(n445) );
  XNOR2_X1 U385 ( .A(n347), .B(n346), .ZN(G51) );
  NAND2_X1 U386 ( .A1(n354), .A2(n353), .ZN(n347) );
  XNOR2_X1 U387 ( .A(n349), .B(n348), .ZN(G57) );
  NAND2_X1 U388 ( .A1(n351), .A2(n350), .ZN(n349) );
  XNOR2_X1 U389 ( .A(n659), .B(n352), .ZN(n351) );
  XNOR2_X1 U390 ( .A(n642), .B(n355), .ZN(n354) );
  INV_X1 U391 ( .A(n641), .ZN(n355) );
  XNOR2_X2 U392 ( .A(n496), .B(n511), .ZN(n657) );
  XNOR2_X2 U393 ( .A(n357), .B(n356), .ZN(n702) );
  NAND2_X1 U394 ( .A1(n561), .A2(n686), .ZN(n357) );
  XNOR2_X2 U395 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n567) );
  XNOR2_X2 U396 ( .A(G902), .B(KEYINPUT15), .ZN(n634) );
  AND2_X2 U397 ( .A1(n375), .A2(KEYINPUT66), .ZN(n374) );
  XNOR2_X1 U398 ( .A(G143), .B(G104), .ZN(n514) );
  XOR2_X1 U399 ( .A(G110), .B(G128), .Z(n467) );
  INV_X1 U400 ( .A(G146), .ZN(n431) );
  NAND2_X2 U401 ( .A1(n393), .A2(n392), .ZN(n388) );
  BUF_X2 U402 ( .A(n556), .Z(n693) );
  NAND2_X1 U403 ( .A1(n414), .A2(n413), .ZN(n392) );
  NOR2_X1 U404 ( .A1(n770), .A2(n771), .ZN(n422) );
  XNOR2_X1 U405 ( .A(n618), .B(KEYINPUT40), .ZN(n770) );
  AND2_X1 U406 ( .A1(n625), .A2(n589), .ZN(n618) );
  AND2_X1 U407 ( .A1(n676), .A2(n706), .ZN(n602) );
  XNOR2_X1 U408 ( .A(n608), .B(n607), .ZN(n707) );
  XNOR2_X1 U409 ( .A(n605), .B(n406), .ZN(n606) );
  XNOR2_X1 U410 ( .A(n639), .B(n640), .ZN(n641) );
  XNOR2_X1 U411 ( .A(n753), .B(n431), .ZN(n511) );
  XNOR2_X1 U412 ( .A(G107), .B(G104), .ZN(n504) );
  XOR2_X2 U413 ( .A(G143), .B(G128), .Z(n531) );
  XNOR2_X1 U414 ( .A(KEYINPUT80), .B(G110), .ZN(n503) );
  XNOR2_X1 U415 ( .A(G116), .B(KEYINPUT77), .ZN(n490) );
  XNOR2_X1 U416 ( .A(KEYINPUT89), .B(KEYINPUT75), .ZN(n489) );
  NAND2_X1 U417 ( .A1(n369), .A2(n444), .ZN(n400) );
  XNOR2_X2 U418 ( .A(n358), .B(KEYINPUT87), .ZN(n591) );
  NAND2_X2 U419 ( .A1(n544), .A2(n703), .ZN(n358) );
  AND2_X1 U420 ( .A1(n369), .A2(n610), .ZN(n676) );
  AND2_X1 U421 ( .A1(n359), .A2(n420), .ZN(n419) );
  XNOR2_X1 U422 ( .A(n602), .B(KEYINPUT47), .ZN(n359) );
  AND2_X1 U423 ( .A1(n421), .A2(n417), .ZN(n619) );
  NAND2_X1 U424 ( .A1(n398), .A2(n397), .ZN(n360) );
  NAND2_X1 U425 ( .A1(n398), .A2(n397), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n379), .B(n367), .ZN(n370) );
  BUF_X1 U427 ( .A(n384), .Z(n361) );
  XNOR2_X2 U428 ( .A(n747), .B(n373), .ZN(n638) );
  XNOR2_X1 U429 ( .A(n486), .B(n432), .ZN(n753) );
  XNOR2_X1 U430 ( .A(n485), .B(G137), .ZN(n433) );
  XOR2_X1 U431 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n465) );
  INV_X1 U432 ( .A(n403), .ZN(n402) );
  INV_X1 U433 ( .A(n604), .ZN(n420) );
  XNOR2_X1 U434 ( .A(n418), .B(KEYINPUT73), .ZN(n417) );
  XNOR2_X1 U435 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n534) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n532) );
  INV_X1 U437 ( .A(n584), .ZN(n415) );
  INV_X1 U438 ( .A(KEYINPUT38), .ZN(n406) );
  XNOR2_X1 U439 ( .A(n380), .B(n495), .ZN(n496) );
  INV_X1 U440 ( .A(G134), .ZN(n454) );
  XNOR2_X1 U441 ( .A(n517), .B(n396), .ZN(n395) );
  INV_X1 U442 ( .A(G122), .ZN(n396) );
  XNOR2_X1 U443 ( .A(G113), .B(G131), .ZN(n517) );
  XNOR2_X1 U444 ( .A(n559), .B(KEYINPUT22), .ZN(n577) );
  NAND2_X1 U445 ( .A1(n578), .A2(n440), .ZN(n439) );
  XNOR2_X1 U446 ( .A(n525), .B(n524), .ZN(n574) );
  INV_X1 U447 ( .A(KEYINPUT86), .ZN(n575) );
  INV_X1 U448 ( .A(G131), .ZN(n485) );
  NAND2_X1 U449 ( .A1(n633), .A2(n368), .ZN(n397) );
  XNOR2_X1 U450 ( .A(KEYINPUT76), .B(G113), .ZN(n487) );
  OR2_X1 U451 ( .A1(n606), .A2(n703), .ZN(n705) );
  NAND2_X1 U452 ( .A1(n606), .A2(n703), .ZN(n608) );
  INV_X1 U453 ( .A(KEYINPUT36), .ZN(n429) );
  INV_X1 U454 ( .A(KEYINPUT34), .ZN(n563) );
  INV_X1 U455 ( .A(G953), .ZN(n441) );
  INV_X1 U456 ( .A(G140), .ZN(n506) );
  INV_X1 U457 ( .A(n606), .ZN(n405) );
  NOR2_X1 U458 ( .A1(n593), .A2(n429), .ZN(n425) );
  XNOR2_X1 U459 ( .A(n516), .B(n395), .ZN(n520) );
  AND2_X1 U460 ( .A1(n643), .A2(G953), .ZN(n737) );
  INV_X2 U461 ( .A(G953), .ZN(n757) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n771) );
  INV_X1 U463 ( .A(KEYINPUT42), .ZN(n407) );
  NAND2_X1 U464 ( .A1(n402), .A2(n401), .ZN(n570) );
  INV_X1 U465 ( .A(n698), .ZN(n401) );
  INV_X1 U466 ( .A(KEYINPUT67), .ZN(n437) );
  AND2_X1 U467 ( .A1(n574), .A2(n565), .ZN(n362) );
  AND2_X1 U468 ( .A1(n755), .A2(n633), .ZN(n363) );
  AND2_X1 U469 ( .A1(n704), .A2(n688), .ZN(n364) );
  INV_X1 U470 ( .A(G146), .ZN(n463) );
  AND2_X1 U471 ( .A1(n706), .A2(n575), .ZN(n365) );
  XOR2_X1 U472 ( .A(n545), .B(KEYINPUT69), .Z(n366) );
  XNOR2_X1 U473 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n367) );
  NAND2_X1 U474 ( .A1(n630), .A2(KEYINPUT68), .ZN(n368) );
  XNOR2_X2 U475 ( .A(n372), .B(n541), .ZN(n544) );
  NAND2_X1 U476 ( .A1(n363), .A2(n370), .ZN(n398) );
  NAND2_X1 U477 ( .A1(n370), .A2(n441), .ZN(n744) );
  XNOR2_X1 U478 ( .A(n371), .B(G119), .ZN(n488) );
  XNOR2_X2 U479 ( .A(G101), .B(KEYINPUT3), .ZN(n371) );
  NAND2_X1 U480 ( .A1(n638), .A2(n634), .ZN(n372) );
  XNOR2_X1 U481 ( .A(n539), .B(n538), .ZN(n373) );
  XNOR2_X2 U482 ( .A(n530), .B(n529), .ZN(n747) );
  NAND2_X1 U483 ( .A1(n376), .A2(n360), .ZN(n637) );
  NAND2_X1 U484 ( .A1(n399), .A2(KEYINPUT2), .ZN(n376) );
  NAND2_X1 U485 ( .A1(n374), .A2(n376), .ZN(n386) );
  XNOR2_X2 U486 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n377) );
  XNOR2_X2 U487 ( .A(G146), .B(G125), .ZN(n378) );
  INV_X1 U488 ( .A(n693), .ZN(n440) );
  NAND2_X1 U489 ( .A1(n389), .A2(n388), .ZN(n379) );
  NAND2_X1 U490 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n579) );
  NOR2_X1 U492 ( .A1(n577), .A2(n439), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n387), .B(n367), .ZN(n629) );
  XNOR2_X1 U494 ( .A(n463), .B(G125), .ZN(n381) );
  XNOR2_X1 U495 ( .A(n484), .B(KEYINPUT4), .ZN(n382) );
  AND2_X1 U496 ( .A1(n436), .A2(n383), .ZN(n414) );
  NOR2_X1 U497 ( .A1(n664), .A2(n575), .ZN(n383) );
  XNOR2_X1 U498 ( .A(n568), .B(n567), .ZN(n384) );
  NAND2_X1 U499 ( .A1(n637), .A2(n636), .ZN(n385) );
  NAND2_X2 U500 ( .A1(n386), .A2(n385), .ZN(n724) );
  INV_X1 U501 ( .A(n664), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n568), .B(n567), .ZN(n663) );
  AND2_X2 U503 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X1 U504 ( .A1(n415), .A2(KEYINPUT44), .ZN(n390) );
  NAND2_X1 U505 ( .A1(n410), .A2(n584), .ZN(n391) );
  INV_X1 U506 ( .A(n394), .ZN(n393) );
  NAND2_X1 U507 ( .A1(n412), .A2(n411), .ZN(n394) );
  XNOR2_X2 U508 ( .A(n492), .B(n491), .ZN(n530) );
  NAND2_X1 U509 ( .A1(n436), .A2(n435), .ZN(n416) );
  NAND2_X1 U510 ( .A1(n620), .A2(n429), .ZN(n428) );
  NAND2_X1 U511 ( .A1(n590), .A2(n596), .ZN(n620) );
  NAND2_X1 U512 ( .A1(n684), .A2(n635), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n629), .A2(n755), .ZN(n684) );
  XNOR2_X2 U514 ( .A(n400), .B(KEYINPUT0), .ZN(n403) );
  NAND2_X1 U515 ( .A1(n402), .A2(n364), .ZN(n559) );
  XNOR2_X1 U516 ( .A(n403), .B(n442), .ZN(n404) );
  XNOR2_X1 U517 ( .A(n381), .B(G140), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n404), .A2(n443), .ZN(n564) );
  NAND2_X1 U519 ( .A1(n404), .A2(n550), .ZN(n551) );
  XNOR2_X1 U520 ( .A(n382), .B(n433), .ZN(n432) );
  NAND2_X1 U521 ( .A1(n716), .A2(n610), .ZN(n408) );
  NAND2_X1 U522 ( .A1(n707), .A2(n704), .ZN(n409) );
  XNOR2_X1 U523 ( .A(n576), .B(KEYINPUT70), .ZN(n410) );
  NAND2_X1 U524 ( .A1(n434), .A2(n365), .ZN(n411) );
  NAND2_X1 U525 ( .A1(n416), .A2(n575), .ZN(n412) );
  NAND2_X1 U526 ( .A1(n434), .A2(n706), .ZN(n413) );
  NOR2_X2 U527 ( .A1(n588), .A2(n577), .ZN(n581) );
  XNOR2_X1 U528 ( .A(n572), .B(KEYINPUT98), .ZN(n434) );
  NAND2_X1 U529 ( .A1(n553), .A2(n440), .ZN(n666) );
  INV_X1 U530 ( .A(n552), .ZN(n553) );
  NAND2_X1 U531 ( .A1(n603), .A2(n419), .ZN(n418) );
  XNOR2_X1 U532 ( .A(n422), .B(KEYINPUT46), .ZN(n421) );
  NAND2_X1 U533 ( .A1(n423), .A2(n425), .ZN(n424) );
  INV_X1 U534 ( .A(n620), .ZN(n423) );
  NAND2_X1 U535 ( .A1(n426), .A2(n424), .ZN(n430) );
  AND2_X1 U536 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U537 ( .A1(n593), .A2(n429), .ZN(n427) );
  NAND2_X1 U538 ( .A1(n430), .A2(n686), .ZN(n594) );
  NAND2_X1 U539 ( .A1(n384), .A2(KEYINPUT44), .ZN(n436) );
  INV_X1 U540 ( .A(KEYINPUT94), .ZN(n442) );
  INV_X1 U541 ( .A(n702), .ZN(n443) );
  BUF_X1 U542 ( .A(n724), .Z(n732) );
  XOR2_X1 U543 ( .A(n549), .B(KEYINPUT93), .Z(n444) );
  INV_X1 U544 ( .A(KEYINPUT85), .ZN(n595) );
  NAND2_X1 U545 ( .A1(n666), .A2(n571), .ZN(n572) );
  XNOR2_X1 U546 ( .A(n507), .B(n506), .ZN(n508) );
  INV_X1 U547 ( .A(KEYINPUT106), .ZN(n607) );
  XNOR2_X1 U548 ( .A(n538), .B(n508), .ZN(n509) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n449) );
  NAND2_X1 U550 ( .A1(n757), .A2(G234), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n447), .B(n446), .ZN(n469) );
  NAND2_X1 U552 ( .A1(G217), .A2(n469), .ZN(n448) );
  XNOR2_X1 U553 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U554 ( .A(KEYINPUT9), .B(G107), .Z(n451) );
  XNOR2_X1 U555 ( .A(G116), .B(G122), .ZN(n450) );
  XNOR2_X1 U556 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U558 ( .A(n531), .B(n454), .ZN(n486) );
  XNOR2_X1 U559 ( .A(n455), .B(n486), .ZN(n646) );
  INV_X1 U560 ( .A(G902), .ZN(n522) );
  NAND2_X1 U561 ( .A1(n646), .A2(n522), .ZN(n458) );
  INV_X1 U562 ( .A(KEYINPUT100), .ZN(n456) );
  XNOR2_X1 U563 ( .A(n456), .B(G478), .ZN(n457) );
  XNOR2_X1 U564 ( .A(n458), .B(n457), .ZN(n573) );
  XOR2_X1 U565 ( .A(KEYINPUT25), .B(KEYINPUT82), .Z(n462) );
  XOR2_X1 U566 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n460) );
  NAND2_X1 U567 ( .A1(G234), .A2(n634), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n460), .B(n459), .ZN(n476) );
  NAND2_X1 U569 ( .A1(n476), .A2(G217), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n475) );
  XNOR2_X1 U571 ( .A(G119), .B(G137), .ZN(n466) );
  XNOR2_X1 U572 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U573 ( .A(n752), .B(n468), .ZN(n473) );
  XOR2_X1 U574 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n471) );
  NAND2_X1 U575 ( .A1(G221), .A2(n469), .ZN(n470) );
  XNOR2_X1 U576 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U577 ( .A(n473), .B(n472), .ZN(n733) );
  XOR2_X1 U578 ( .A(n475), .B(n474), .Z(n587) );
  NAND2_X1 U579 ( .A1(n476), .A2(G221), .ZN(n477) );
  XOR2_X1 U580 ( .A(KEYINPUT21), .B(n477), .Z(n688) );
  NAND2_X1 U581 ( .A1(G234), .A2(G237), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n478), .B(KEYINPUT14), .ZN(n480) );
  NAND2_X1 U583 ( .A1(G952), .A2(n480), .ZN(n715) );
  NOR2_X1 U584 ( .A1(n715), .A2(G953), .ZN(n479) );
  XNOR2_X1 U585 ( .A(n479), .B(KEYINPUT91), .ZN(n548) );
  NAND2_X1 U586 ( .A1(G902), .A2(n480), .ZN(n546) );
  NOR2_X1 U587 ( .A1(G900), .A2(n546), .ZN(n481) );
  NAND2_X1 U588 ( .A1(G953), .A2(n481), .ZN(n482) );
  NAND2_X1 U589 ( .A1(n548), .A2(n482), .ZN(n613) );
  NAND2_X1 U590 ( .A1(n445), .A2(n613), .ZN(n483) );
  NOR2_X1 U591 ( .A1(n573), .A2(n483), .ZN(n528) );
  XOR2_X1 U592 ( .A(KEYINPUT103), .B(KEYINPUT30), .Z(n502) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U595 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n494) );
  NOR2_X1 U596 ( .A1(G953), .A2(G237), .ZN(n518) );
  NAND2_X1 U597 ( .A1(n518), .A2(G210), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U599 ( .A1(n657), .A2(n522), .ZN(n499) );
  INV_X1 U600 ( .A(KEYINPUT97), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n497), .B(G472), .ZN(n498) );
  XNOR2_X2 U602 ( .A(n499), .B(n498), .ZN(n556) );
  INV_X1 U603 ( .A(G237), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n522), .A2(n500), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n556), .A2(n703), .ZN(n501) );
  XNOR2_X1 U606 ( .A(n502), .B(n501), .ZN(n612) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n746) );
  XNOR2_X1 U608 ( .A(n746), .B(KEYINPUT78), .ZN(n538) );
  NAND2_X1 U609 ( .A1(G227), .A2(n757), .ZN(n505) );
  XOR2_X1 U610 ( .A(n505), .B(KEYINPUT83), .Z(n507) );
  XNOR2_X1 U611 ( .A(n509), .B(G101), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n511), .B(n510), .ZN(n728) );
  NOR2_X1 U613 ( .A1(G902), .A2(n728), .ZN(n513) );
  INV_X1 U614 ( .A(G469), .ZN(n512) );
  XNOR2_X2 U615 ( .A(n513), .B(n512), .ZN(n599) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n515) );
  XNOR2_X1 U617 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U618 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U620 ( .A(n521), .B(n752), .ZN(n652) );
  NAND2_X1 U621 ( .A1(n652), .A2(n522), .ZN(n525) );
  INV_X1 U622 ( .A(KEYINPUT13), .ZN(n523) );
  XNOR2_X1 U623 ( .A(n523), .B(G475), .ZN(n524) );
  NAND2_X1 U624 ( .A1(n599), .A2(n574), .ZN(n526) );
  NOR2_X1 U625 ( .A1(n612), .A2(n526), .ZN(n527) );
  NAND2_X1 U626 ( .A1(n528), .A2(n527), .ZN(n543) );
  XNOR2_X1 U627 ( .A(KEYINPUT16), .B(G122), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n532), .B(n531), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n757), .A2(G224), .ZN(n533) );
  XNOR2_X1 U630 ( .A(n533), .B(KEYINPUT18), .ZN(n535) );
  XNOR2_X1 U631 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n537), .B(n536), .ZN(n539) );
  AND2_X1 U633 ( .A1(n540), .A2(G210), .ZN(n541) );
  BUF_X1 U634 ( .A(n544), .Z(n605) );
  INV_X1 U635 ( .A(n605), .ZN(n542) );
  NOR2_X1 U636 ( .A1(n543), .A2(n542), .ZN(n604) );
  XOR2_X1 U637 ( .A(G143), .B(n604), .Z(G45) );
  XNOR2_X1 U638 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n545) );
  XNOR2_X1 U639 ( .A(G898), .B(KEYINPUT92), .ZN(n741) );
  OR2_X1 U640 ( .A1(n757), .A2(n741), .ZN(n748) );
  OR2_X1 U641 ( .A1(n546), .A2(n748), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U643 ( .A1(n599), .A2(n445), .ZN(n611) );
  INV_X1 U644 ( .A(n611), .ZN(n550) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT96), .ZN(n552) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n617) );
  NOR2_X1 U647 ( .A1(n666), .A2(n617), .ZN(n554) );
  XOR2_X1 U648 ( .A(G104), .B(n554), .Z(G6) );
  INV_X1 U649 ( .A(KEYINPUT6), .ZN(n555) );
  XNOR2_X1 U650 ( .A(n556), .B(n555), .ZN(n588) );
  INV_X1 U651 ( .A(n574), .ZN(n557) );
  NAND2_X1 U652 ( .A1(n573), .A2(n557), .ZN(n558) );
  XNOR2_X1 U653 ( .A(KEYINPUT101), .B(n558), .ZN(n704) );
  XNOR2_X2 U654 ( .A(n599), .B(KEYINPUT1), .ZN(n686) );
  INV_X1 U655 ( .A(n587), .ZN(n689) );
  NOR2_X1 U656 ( .A1(n686), .A2(n689), .ZN(n560) );
  AND2_X1 U657 ( .A1(n581), .A2(n560), .ZN(n664) );
  AND2_X1 U658 ( .A1(n588), .A2(n445), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n564), .B(n563), .ZN(n566) );
  INV_X1 U660 ( .A(n573), .ZN(n565) );
  NAND2_X1 U661 ( .A1(n566), .A2(n362), .ZN(n568) );
  AND2_X1 U662 ( .A1(n686), .A2(n445), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n569), .A2(n693), .ZN(n698) );
  XNOR2_X1 U664 ( .A(n570), .B(KEYINPUT31), .ZN(n681) );
  INV_X1 U665 ( .A(n681), .ZN(n571) );
  OR2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n665) );
  NAND2_X1 U667 ( .A1(n617), .A2(n665), .ZN(n706) );
  NOR2_X2 U668 ( .A1(n663), .A2(KEYINPUT44), .ZN(n576) );
  INV_X1 U669 ( .A(n686), .ZN(n578) );
  AND2_X1 U670 ( .A1(n579), .A2(n689), .ZN(n671) );
  AND2_X1 U671 ( .A1(n686), .A2(n689), .ZN(n580) );
  NAND2_X1 U672 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U673 ( .A(KEYINPUT32), .ZN(n582) );
  XNOR2_X1 U674 ( .A(n583), .B(n582), .ZN(n769) );
  NOR2_X2 U675 ( .A1(n671), .A2(n769), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n688), .A2(n613), .ZN(n585) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n585), .ZN(n586) );
  NOR2_X1 U678 ( .A1(n587), .A2(n586), .ZN(n596) );
  INV_X1 U679 ( .A(n617), .ZN(n589) );
  AND2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n590) );
  BUF_X1 U681 ( .A(n591), .Z(n592) );
  INV_X1 U682 ( .A(n592), .ZN(n593) );
  XNOR2_X1 U683 ( .A(n594), .B(KEYINPUT108), .ZN(n767) );
  XNOR2_X1 U684 ( .A(n767), .B(n595), .ZN(n603) );
  XOR2_X1 U685 ( .A(KEYINPUT104), .B(KEYINPUT28), .Z(n598) );
  NAND2_X1 U686 ( .A1(n693), .A2(n596), .ZN(n597) );
  XNOR2_X1 U687 ( .A(n598), .B(n597), .ZN(n600) );
  NAND2_X1 U688 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U689 ( .A(n601), .B(KEYINPUT105), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n609) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U693 ( .A(n616), .B(KEYINPUT39), .Z(n625) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT48), .ZN(n628) );
  NOR2_X1 U695 ( .A1(n620), .A2(n686), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n621), .A2(n703), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT43), .B(n622), .Z(n623) );
  NOR2_X1 U698 ( .A1(n623), .A2(n605), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT102), .ZN(n766) );
  INV_X1 U700 ( .A(n665), .ZN(n680) );
  NAND2_X1 U701 ( .A1(n625), .A2(n680), .ZN(n683) );
  INV_X1 U702 ( .A(n683), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n766), .A2(n626), .ZN(n627) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT68), .ZN(n632) );
  INV_X1 U706 ( .A(n634), .ZN(n631) );
  OR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U708 ( .A1(n634), .A2(KEYINPUT68), .ZN(n635) );
  INV_X1 U709 ( .A(KEYINPUT66), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n724), .A2(G210), .ZN(n642) );
  BUF_X1 U711 ( .A(n638), .Z(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n640) );
  INV_X1 U713 ( .A(G952), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n724), .A2(G478), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X2 U716 ( .A1(n649), .A2(n737), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT120), .ZN(G63) );
  NAND2_X1 U718 ( .A1(n724), .A2(G475), .ZN(n654) );
  XNOR2_X1 U719 ( .A(KEYINPUT118), .B(KEYINPUT59), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U721 ( .A1(n655), .A2(n737), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n656), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U723 ( .A1(n724), .A2(G472), .ZN(n659) );
  XOR2_X1 U724 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n661) );
  XOR2_X1 U725 ( .A(n361), .B(G122), .Z(G24) );
  XOR2_X1 U726 ( .A(G101), .B(n664), .Z(G3) );
  XOR2_X1 U727 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n668) );
  NOR2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U729 ( .A(n668), .B(n667), .Z(n670) );
  XOR2_X1 U730 ( .A(G107), .B(KEYINPUT26), .Z(n669) );
  XNOR2_X1 U731 ( .A(n670), .B(n669), .ZN(G9) );
  XOR2_X1 U732 ( .A(G110), .B(n671), .Z(n672) );
  XNOR2_X1 U733 ( .A(KEYINPUT110), .B(n672), .ZN(G12) );
  AND2_X1 U734 ( .A1(n676), .A2(n680), .ZN(n674) );
  XNOR2_X1 U735 ( .A(KEYINPUT111), .B(KEYINPUT29), .ZN(n673) );
  XNOR2_X1 U736 ( .A(n674), .B(n673), .ZN(n675) );
  XOR2_X1 U737 ( .A(G128), .B(n675), .Z(G30) );
  AND2_X1 U738 ( .A1(n676), .A2(n589), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT112), .B(n677), .Z(n678) );
  XNOR2_X1 U740 ( .A(G146), .B(n678), .ZN(G48) );
  NAND2_X1 U741 ( .A1(n681), .A2(n589), .ZN(n679) );
  XNOR2_X1 U742 ( .A(n679), .B(G113), .ZN(G15) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U744 ( .A(n682), .B(G116), .ZN(G18) );
  XNOR2_X1 U745 ( .A(G134), .B(n683), .ZN(G36) );
  BUF_X1 U746 ( .A(n684), .Z(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT2), .ZN(n721) );
  NOR2_X1 U748 ( .A1(n445), .A2(n686), .ZN(n687) );
  XOR2_X1 U749 ( .A(KEYINPUT50), .B(n687), .Z(n696) );
  XOR2_X1 U750 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n692) );
  INV_X1 U751 ( .A(n688), .ZN(n690) );
  NAND2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U753 ( .A(n692), .B(n691), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n699) );
  XNOR2_X1 U758 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U759 ( .A1(n716), .A2(n701), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U761 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n443), .A2(n710), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U765 ( .A(KEYINPUT52), .B(n713), .Z(n714) );
  NOR2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n718) );
  AND2_X1 U767 ( .A1(n443), .A2(n716), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT115), .B(n719), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n757), .A2(n722), .ZN(n723) );
  XOR2_X1 U772 ( .A(KEYINPUT53), .B(n723), .Z(G75) );
  NAND2_X1 U773 ( .A1(n732), .A2(G469), .ZN(n730) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n726) );
  XNOR2_X1 U775 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n727) );
  XOR2_X1 U777 ( .A(n728), .B(n727), .Z(n729) );
  XNOR2_X1 U778 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n737), .A2(n731), .ZN(G54) );
  NAND2_X1 U780 ( .A1(n732), .A2(G217), .ZN(n735) );
  XOR2_X1 U781 ( .A(n733), .B(KEYINPUT121), .Z(n734) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U783 ( .A1(n737), .A2(n736), .ZN(G66) );
  XOR2_X1 U784 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n739) );
  NAND2_X1 U785 ( .A1(G224), .A2(G953), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(KEYINPUT122), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U790 ( .A(n745), .B(KEYINPUT124), .ZN(n751) );
  XNOR2_X1 U791 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U792 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U793 ( .A(n751), .B(n750), .Z(G69) );
  XOR2_X1 U794 ( .A(n753), .B(n752), .Z(n754) );
  XNOR2_X1 U795 ( .A(KEYINPUT125), .B(n754), .ZN(n760) );
  INV_X1 U796 ( .A(n760), .ZN(n756) );
  XNOR2_X1 U797 ( .A(n756), .B(n755), .ZN(n758) );
  NAND2_X1 U798 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n759), .ZN(n765) );
  XNOR2_X1 U800 ( .A(G227), .B(n760), .ZN(n761) );
  NAND2_X1 U801 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U802 ( .A1(G953), .A2(n762), .ZN(n763) );
  XOR2_X1 U803 ( .A(KEYINPUT127), .B(n763), .Z(n764) );
  NAND2_X1 U804 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U805 ( .A(G140), .B(n766), .Z(G42) );
  XOR2_X1 U806 ( .A(G125), .B(n767), .Z(n768) );
  XNOR2_X1 U807 ( .A(KEYINPUT37), .B(n768), .ZN(G27) );
  XOR2_X1 U808 ( .A(G119), .B(n769), .Z(G21) );
  XOR2_X1 U809 ( .A(G131), .B(n770), .Z(G33) );
  XOR2_X1 U810 ( .A(n771), .B(G137), .Z(G39) );
endmodule

