

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n583), .A2(n582), .ZN(G164) );
  INV_X1 U556 ( .A(n672), .ZN(n658) );
  XNOR2_X1 U557 ( .A(KEYINPUT65), .B(n557), .ZN(n801) );
  XNOR2_X1 U558 ( .A(n681), .B(KEYINPUT32), .ZN(n700) );
  XNOR2_X1 U559 ( .A(n628), .B(n536), .ZN(n648) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n536) );
  AND2_X1 U561 ( .A1(n689), .A2(n704), .ZN(n690) );
  NAND2_X1 U562 ( .A1(n730), .A2(n625), .ZN(n672) );
  INV_X1 U563 ( .A(KEYINPUT99), .ZN(n678) );
  OR2_X1 U564 ( .A1(n648), .A2(n962), .ZN(n647) );
  NOR2_X1 U565 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U566 ( .A(n526), .B(n525), .ZN(n524) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n525) );
  AND2_X1 U568 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U569 ( .A1(n521), .A2(n535), .ZN(n534) );
  AND2_X1 U570 ( .A1(n957), .A2(n523), .ZN(n533) );
  XNOR2_X1 U571 ( .A(n530), .B(n707), .ZN(n529) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n730) );
  XNOR2_X1 U573 ( .A(n537), .B(n576), .ZN(n577) );
  INV_X1 U574 ( .A(KEYINPUT89), .ZN(n576) );
  OR2_X1 U575 ( .A1(G2105), .A2(n541), .ZN(n542) );
  AND2_X1 U576 ( .A1(n695), .A2(n694), .ZN(n521) );
  XNOR2_X1 U577 ( .A(KEYINPUT28), .B(n657), .ZN(n522) );
  OR2_X1 U578 ( .A1(n710), .A2(n697), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n662), .ZN(n671) );
  NAND2_X1 U580 ( .A1(n527), .A2(n522), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n655), .B(n528), .ZN(n527) );
  INV_X1 U582 ( .A(KEYINPUT97), .ZN(n528) );
  NOR2_X1 U583 ( .A1(n531), .A2(n529), .ZN(n745) );
  NAND2_X1 U584 ( .A1(n706), .A2(n705), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n532), .A2(n712), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n532) );
  INV_X1 U587 ( .A(KEYINPUT33), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n901), .A2(G138), .ZN(n537) );
  XNOR2_X2 U589 ( .A(n538), .B(KEYINPUT17), .ZN(n901) );
  NAND2_X1 U590 ( .A1(n579), .A2(n546), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT27), .B(n649), .Z(n539) );
  AND2_X1 U592 ( .A1(n644), .A2(n643), .ZN(n540) );
  AND2_X1 U593 ( .A1(n645), .A2(n540), .ZN(n646) );
  NOR2_X1 U594 ( .A1(n555), .A2(G651), .ZN(n797) );
  NOR2_X1 U595 ( .A1(G543), .A2(G651), .ZN(n794) );
  XOR2_X1 U596 ( .A(n624), .B(n623), .Z(n962) );
  NOR2_X1 U597 ( .A1(n550), .A2(n549), .ZN(G160) );
  NAND2_X1 U598 ( .A1(G2104), .A2(G101), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT64), .B(n542), .Z(n543) );
  XNOR2_X1 U600 ( .A(n543), .B(KEYINPUT23), .ZN(n545) );
  INV_X1 U601 ( .A(G2104), .ZN(n579) );
  INV_X1 U602 ( .A(G2105), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n579), .A2(n546), .ZN(n905) );
  NAND2_X1 U604 ( .A1(G113), .A2(n905), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n901), .A2(G137), .ZN(n548) );
  NOR2_X1 U607 ( .A1(G2104), .A2(n546), .ZN(n906) );
  NAND2_X1 U608 ( .A1(G125), .A2(n906), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U610 ( .A(KEYINPUT0), .B(G543), .Z(n555) );
  NAND2_X1 U611 ( .A1(n797), .A2(G48), .ZN(n562) );
  INV_X1 U612 ( .A(G651), .ZN(n556) );
  NOR2_X1 U613 ( .A1(G543), .A2(n556), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT1), .B(n551), .Z(n793) );
  NAND2_X1 U615 ( .A1(G61), .A2(n793), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G86), .A2(n794), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT82), .B(n554), .ZN(n560) );
  OR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n801), .A2(G73), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT2), .B(n558), .Z(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT83), .B(n563), .Z(G305) );
  NAND2_X1 U625 ( .A1(n794), .A2(G89), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G76), .A2(n801), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n567), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n797), .A2(G51), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT71), .B(n568), .Z(n570) );
  NAND2_X1 U632 ( .A1(n793), .A2(G63), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT6), .B(n571), .Z(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U636 ( .A(KEYINPUT7), .B(n574), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT72), .B(n575), .ZN(G286) );
  NAND2_X1 U639 ( .A1(n905), .A2(G114), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n583) );
  NOR2_X1 U641 ( .A1(G2105), .A2(n579), .ZN(n902) );
  NAND2_X1 U642 ( .A1(G102), .A2(n902), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G126), .A2(n906), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G65), .A2(n793), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G53), .A2(n797), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(n586), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G91), .A2(n794), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G78), .A2(n801), .ZN(n587) );
  AND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(G299) );
  NAND2_X1 U653 ( .A1(G64), .A2(n793), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G52), .A2(n797), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n597) );
  NAND2_X1 U656 ( .A1(G90), .A2(n794), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G77), .A2(n801), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT9), .B(n595), .Z(n596) );
  NOR2_X1 U660 ( .A1(n597), .A2(n596), .ZN(G171) );
  NAND2_X1 U661 ( .A1(G50), .A2(n797), .ZN(n598) );
  XNOR2_X1 U662 ( .A(n598), .B(KEYINPUT84), .ZN(n600) );
  NAND2_X1 U663 ( .A1(n793), .A2(G62), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U665 ( .A1(G88), .A2(n794), .ZN(n602) );
  NAND2_X1 U666 ( .A1(G75), .A2(n801), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(G166) );
  INV_X1 U669 ( .A(G166), .ZN(G303) );
  NAND2_X1 U670 ( .A1(n555), .A2(G87), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G49), .A2(n797), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G74), .A2(G651), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U674 ( .A1(n793), .A2(n607), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U676 ( .A(KEYINPUT81), .B(n610), .Z(G288) );
  AND2_X1 U677 ( .A1(n794), .A2(G85), .ZN(n614) );
  NAND2_X1 U678 ( .A1(G60), .A2(n793), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G47), .A2(n797), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n801), .A2(G72), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n616), .A2(n615), .ZN(G290) );
  XOR2_X1 U684 ( .A(G1981), .B(G305), .Z(n957) );
  NAND2_X1 U685 ( .A1(G66), .A2(n793), .ZN(n618) );
  NAND2_X1 U686 ( .A1(G92), .A2(n794), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U688 ( .A1(G79), .A2(n801), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G54), .A2(n797), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n624) );
  XNOR2_X1 U692 ( .A(KEYINPUT70), .B(KEYINPUT15), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G160), .A2(G40), .ZN(n729) );
  INV_X1 U694 ( .A(n729), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n658), .A2(G2067), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G1348), .A2(n672), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U698 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n641) );
  NOR2_X1 U699 ( .A1(G1996), .A2(n641), .ZN(n639) );
  XOR2_X1 U700 ( .A(KEYINPUT14), .B(KEYINPUT68), .Z(n630) );
  NAND2_X1 U701 ( .A1(G56), .A2(n793), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n794), .A2(G81), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT12), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G68), .A2(n801), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U707 ( .A(KEYINPUT13), .B(n634), .Z(n635) );
  NOR2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n797), .A2(G43), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n955) );
  NOR2_X1 U711 ( .A1(n639), .A2(n955), .ZN(n645) );
  INV_X1 U712 ( .A(G1341), .ZN(n956) );
  NAND2_X1 U713 ( .A1(n956), .A2(n641), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n640), .A2(n672), .ZN(n644) );
  AND2_X1 U715 ( .A1(G1996), .A2(n658), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n654) );
  AND2_X1 U718 ( .A1(n962), .A2(n648), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n658), .A2(G2072), .ZN(n649) );
  XNOR2_X1 U720 ( .A(G1956), .B(KEYINPUT94), .ZN(n935) );
  NAND2_X1 U721 ( .A1(n672), .A2(n935), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n539), .A2(n650), .ZN(n656) );
  NOR2_X1 U723 ( .A1(n656), .A2(G299), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U725 ( .A1(G299), .A2(n656), .ZN(n657) );
  INV_X1 U726 ( .A(G1961), .ZN(n945) );
  NAND2_X1 U727 ( .A1(n672), .A2(n945), .ZN(n660) );
  XNOR2_X1 U728 ( .A(G2078), .B(KEYINPUT25), .ZN(n1022) );
  NAND2_X1 U729 ( .A1(n658), .A2(n1022), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n666) );
  AND2_X1 U731 ( .A1(n666), .A2(G171), .ZN(n661) );
  XNOR2_X1 U732 ( .A(KEYINPUT93), .B(n661), .ZN(n662) );
  NOR2_X1 U733 ( .A1(G2084), .A2(n672), .ZN(n686) );
  NAND2_X1 U734 ( .A1(G8), .A2(n672), .ZN(n710) );
  NOR2_X1 U735 ( .A1(G1966), .A2(n710), .ZN(n682) );
  NOR2_X1 U736 ( .A1(n686), .A2(n682), .ZN(n663) );
  NAND2_X1 U737 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U738 ( .A(KEYINPUT30), .B(n664), .ZN(n665) );
  NOR2_X1 U739 ( .A1(G168), .A2(n665), .ZN(n668) );
  NOR2_X1 U740 ( .A1(G171), .A2(n666), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT31), .B(n669), .Z(n670) );
  NAND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n684) );
  NAND2_X1 U744 ( .A1(G286), .A2(n684), .ZN(n677) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n710), .ZN(n674) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n675), .A2(G303), .ZN(n676) );
  NAND2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n680), .A2(G8), .ZN(n681) );
  INV_X1 U752 ( .A(n682), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT98), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n686), .A2(G8), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n698) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n969) );
  AND2_X1 U757 ( .A1(n698), .A2(n969), .ZN(n689) );
  INV_X1 U758 ( .A(n710), .ZN(n704) );
  NAND2_X1 U759 ( .A1(n700), .A2(n690), .ZN(n695) );
  INV_X1 U760 ( .A(n969), .ZN(n692) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n696) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n696), .A2(n691), .ZN(n973) );
  OR2_X1 U764 ( .A1(n692), .A2(n973), .ZN(n693) );
  OR2_X1 U765 ( .A1(n710), .A2(n693), .ZN(n694) );
  NAND2_X1 U766 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  AND2_X1 U767 ( .A1(n698), .A2(n710), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n706) );
  NOR2_X1 U769 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U770 ( .A1(G8), .A2(n701), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n702), .B(KEYINPUT100), .ZN(n703) );
  OR2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  INV_X1 U773 ( .A(KEYINPUT101), .ZN(n707) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n708) );
  XOR2_X1 U775 ( .A(n708), .B(KEYINPUT24), .Z(n709) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U777 ( .A(n711), .B(KEYINPUT92), .Z(n712) );
  NAND2_X1 U778 ( .A1(G131), .A2(n901), .ZN(n714) );
  NAND2_X1 U779 ( .A1(G95), .A2(n902), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G107), .A2(n905), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G119), .A2(n906), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n883) );
  INV_X1 U785 ( .A(G1991), .ZN(n1016) );
  NOR2_X1 U786 ( .A1(n883), .A2(n1016), .ZN(n728) );
  NAND2_X1 U787 ( .A1(G141), .A2(n901), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G117), .A2(n905), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U790 ( .A1(G105), .A2(n902), .ZN(n721) );
  XNOR2_X1 U791 ( .A(n721), .B(KEYINPUT38), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n722), .B(KEYINPUT91), .ZN(n723) );
  NOR2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n906), .A2(G129), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n897) );
  AND2_X1 U796 ( .A1(n897), .A2(G1996), .ZN(n727) );
  NOR2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n1003) );
  NOR2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n761) );
  INV_X1 U799 ( .A(n761), .ZN(n731) );
  NOR2_X1 U800 ( .A1(n1003), .A2(n731), .ZN(n752) );
  INV_X1 U801 ( .A(n752), .ZN(n743) );
  XNOR2_X1 U802 ( .A(KEYINPUT37), .B(G2067), .ZN(n759) );
  NAND2_X1 U803 ( .A1(G140), .A2(n901), .ZN(n733) );
  NAND2_X1 U804 ( .A1(G104), .A2(n902), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U806 ( .A(KEYINPUT34), .B(n734), .ZN(n740) );
  NAND2_X1 U807 ( .A1(G116), .A2(n905), .ZN(n736) );
  NAND2_X1 U808 ( .A1(G128), .A2(n906), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U810 ( .A(KEYINPUT35), .B(n737), .Z(n738) );
  XNOR2_X1 U811 ( .A(KEYINPUT90), .B(n738), .ZN(n739) );
  NOR2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n741), .ZN(n916) );
  NOR2_X1 U814 ( .A1(n759), .A2(n916), .ZN(n757) );
  NAND2_X1 U815 ( .A1(n761), .A2(n757), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U818 ( .A(n746), .B(KEYINPUT102), .ZN(n748) );
  XNOR2_X1 U819 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U820 ( .A1(n975), .A2(n761), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n764) );
  XOR2_X1 U822 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n756) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n897), .ZN(n749) );
  XOR2_X1 U824 ( .A(KEYINPUT103), .B(n749), .Z(n992) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n750) );
  AND2_X1 U826 ( .A1(n1016), .A2(n883), .ZN(n999) );
  NOR2_X1 U827 ( .A1(n750), .A2(n999), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n753), .B(KEYINPUT104), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n992), .A2(n754), .ZN(n755) );
  XNOR2_X1 U831 ( .A(n756), .B(n755), .ZN(n758) );
  INV_X1 U832 ( .A(n757), .ZN(n1002) );
  NAND2_X1 U833 ( .A1(n758), .A2(n1002), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n759), .A2(n916), .ZN(n988) );
  NAND2_X1 U835 ( .A1(n760), .A2(n988), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  NAND2_X1 U840 ( .A1(G94), .A2(G452), .ZN(n766) );
  XOR2_X1 U841 ( .A(KEYINPUT66), .B(n766), .Z(G173) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n847) );
  NAND2_X1 U845 ( .A1(n847), .A2(G567), .ZN(n768) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n768), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n774) );
  OR2_X1 U848 ( .A1(n955), .A2(n774), .ZN(G153) );
  INV_X1 U849 ( .A(G868), .ZN(n818) );
  NOR2_X1 U850 ( .A1(n818), .A2(G171), .ZN(n769) );
  XNOR2_X1 U851 ( .A(n769), .B(KEYINPUT69), .ZN(n771) );
  OR2_X1 U852 ( .A1(G868), .A2(n962), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n771), .A2(n770), .ZN(G284) );
  NAND2_X1 U854 ( .A1(G868), .A2(G286), .ZN(n773) );
  NAND2_X1 U855 ( .A1(G299), .A2(n818), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n775), .A2(n962), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n955), .ZN(n777) );
  XOR2_X1 U861 ( .A(KEYINPUT73), .B(n777), .Z(n780) );
  NAND2_X1 U862 ( .A1(G868), .A2(n962), .ZN(n778) );
  NOR2_X1 U863 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G123), .A2(n906), .ZN(n781) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n781), .Z(n787) );
  NAND2_X1 U867 ( .A1(n905), .A2(G111), .ZN(n782) );
  XNOR2_X1 U868 ( .A(n782), .B(KEYINPUT74), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G99), .A2(n902), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U871 ( .A(KEYINPUT75), .B(n785), .Z(n786) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n901), .A2(G135), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n1000) );
  XOR2_X1 U875 ( .A(G2096), .B(KEYINPUT76), .Z(n790) );
  XNOR2_X1 U876 ( .A(n1000), .B(n790), .ZN(n792) );
  INV_X1 U877 ( .A(G2100), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(G156) );
  NAND2_X1 U879 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G93), .A2(n794), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G55), .A2(n797), .ZN(n798) );
  XNOR2_X1 U883 ( .A(KEYINPUT79), .B(n798), .ZN(n799) );
  NOR2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U885 ( .A1(n801), .A2(G80), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n803), .A2(n802), .ZN(n817) );
  NAND2_X1 U887 ( .A1(n962), .A2(G559), .ZN(n804) );
  XOR2_X1 U888 ( .A(n955), .B(n804), .Z(n815) );
  XNOR2_X1 U889 ( .A(KEYINPUT77), .B(n815), .ZN(n805) );
  NOR2_X1 U890 ( .A1(G860), .A2(n805), .ZN(n806) );
  XOR2_X1 U891 ( .A(n806), .B(KEYINPUT78), .Z(n807) );
  XNOR2_X1 U892 ( .A(KEYINPUT80), .B(n807), .ZN(n808) );
  XNOR2_X1 U893 ( .A(n817), .B(n808), .ZN(G145) );
  XOR2_X1 U894 ( .A(G305), .B(G299), .Z(n809) );
  XNOR2_X1 U895 ( .A(n817), .B(n809), .ZN(n810) );
  XNOR2_X1 U896 ( .A(KEYINPUT85), .B(n810), .ZN(n812) );
  XNOR2_X1 U897 ( .A(G290), .B(KEYINPUT19), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U899 ( .A(n813), .B(G288), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n814), .B(G303), .ZN(n871) );
  XNOR2_X1 U901 ( .A(n815), .B(n871), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n816), .A2(G868), .ZN(n820) );
  NAND2_X1 U903 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n821) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n821), .Z(n822) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n822), .ZN(n823) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n823), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n824), .A2(G2072), .ZN(n825) );
  XNOR2_X1 U910 ( .A(KEYINPUT86), .B(n825), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n826) );
  NOR2_X1 U913 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(G108), .A2(n827), .ZN(n852) );
  NAND2_X1 U915 ( .A1(G567), .A2(n852), .ZN(n834) );
  XOR2_X1 U916 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n829) );
  NAND2_X1 U917 ( .A1(G132), .A2(G82), .ZN(n828) );
  XNOR2_X1 U918 ( .A(n829), .B(n828), .ZN(n830) );
  NOR2_X1 U919 ( .A1(n830), .A2(G218), .ZN(n831) );
  XNOR2_X1 U920 ( .A(KEYINPUT88), .B(n831), .ZN(n832) );
  NAND2_X1 U921 ( .A1(n832), .A2(G96), .ZN(n851) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n851), .ZN(n833) );
  NAND2_X1 U923 ( .A1(n834), .A2(n833), .ZN(n853) );
  NAND2_X1 U924 ( .A1(G483), .A2(G661), .ZN(n835) );
  NOR2_X1 U925 ( .A1(n853), .A2(n835), .ZN(n850) );
  NAND2_X1 U926 ( .A1(n850), .A2(G36), .ZN(G176) );
  XNOR2_X1 U927 ( .A(G2443), .B(G2454), .ZN(n845) );
  XOR2_X1 U928 ( .A(KEYINPUT106), .B(G2430), .Z(n837) );
  XNOR2_X1 U929 ( .A(G2446), .B(KEYINPUT107), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U931 ( .A(G2451), .B(G2427), .Z(n839) );
  XNOR2_X1 U932 ( .A(G1348), .B(G1341), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U935 ( .A(G2438), .B(G2435), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U937 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U938 ( .A1(n846), .A2(G14), .ZN(n920) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(n920), .Z(G401) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n847), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U942 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(G188) );
  NOR2_X1 U945 ( .A1(n852), .A2(n851), .ZN(G325) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U948 ( .A(G132), .ZN(G219) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G82), .ZN(G220) );
  INV_X1 U952 ( .A(G69), .ZN(G235) );
  INV_X1 U953 ( .A(n853), .ZN(G319) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1961), .B(G1971), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1976), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(n864), .B(G2474), .Z(n866) );
  XNOR2_X1 U967 ( .A(G1981), .B(G1966), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT41), .B(G1956), .Z(n868) );
  XNOR2_X1 U970 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(G229) );
  INV_X1 U973 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U974 ( .A(G286), .B(n871), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n962), .B(G301), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(n874), .B(n955), .Z(n875) );
  NOR2_X1 U978 ( .A1(G37), .A2(n875), .ZN(G397) );
  NAND2_X1 U979 ( .A1(G124), .A2(n906), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n905), .A2(G112), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G136), .A2(n901), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G100), .A2(n902), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U986 ( .A1(n882), .A2(n881), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n885) );
  XNOR2_X1 U988 ( .A(n883), .B(KEYINPUT113), .ZN(n884) );
  XNOR2_X1 U989 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U990 ( .A(G164), .B(n886), .ZN(n915) );
  XNOR2_X1 U991 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G142), .A2(n901), .ZN(n888) );
  NAND2_X1 U993 ( .A1(G106), .A2(n902), .ZN(n887) );
  NAND2_X1 U994 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U995 ( .A(n889), .B(KEYINPUT45), .ZN(n890) );
  XNOR2_X1 U996 ( .A(n891), .B(n890), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n906), .A2(G130), .ZN(n892) );
  XNOR2_X1 U998 ( .A(n892), .B(KEYINPUT110), .ZN(n894) );
  NAND2_X1 U999 ( .A1(G118), .A2(n905), .ZN(n893) );
  NAND2_X1 U1000 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U1001 ( .A1(n896), .A2(n895), .ZN(n899) );
  XOR2_X1 U1002 ( .A(G162), .B(n897), .Z(n898) );
  XNOR2_X1 U1003 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1004 ( .A(n1000), .B(n900), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n901), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n902), .ZN(n903) );
  NAND2_X1 U1007 ( .A1(n904), .A2(n903), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n905), .ZN(n908) );
  NAND2_X1 U1009 ( .A1(G127), .A2(n906), .ZN(n907) );
  NAND2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1011 ( .A(KEYINPUT47), .B(n909), .Z(n910) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n984) );
  XNOR2_X1 U1013 ( .A(G160), .B(n984), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1016 ( .A(n917), .B(n916), .Z(n918) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n918), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT114), .B(n919), .ZN(G395) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n920), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n921), .Z(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(KEYINPUT115), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT116), .B(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(G397), .A2(G395), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1029 ( .A(G1976), .B(G23), .Z(n929) );
  XOR2_X1 U1030 ( .A(G1971), .B(G22), .Z(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G24), .B(G1986), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1034 ( .A(KEYINPUT58), .B(n932), .Z(n952) );
  XOR2_X1 U1035 ( .A(KEYINPUT126), .B(G4), .Z(n934) );
  XNOR2_X1 U1036 ( .A(G1348), .B(KEYINPUT59), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(n934), .B(n933), .ZN(n943) );
  XOR2_X1 U1038 ( .A(n935), .B(G20), .Z(n940) );
  XNOR2_X1 U1039 ( .A(G1981), .B(G6), .ZN(n937) );
  XNOR2_X1 U1040 ( .A(G19), .B(G1341), .ZN(n936) );
  NOR2_X1 U1041 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1042 ( .A(n938), .B(KEYINPUT124), .ZN(n939) );
  NAND2_X1 U1043 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1044 ( .A(KEYINPUT125), .B(n941), .Z(n942) );
  NOR2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT60), .B(n944), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n945), .B(G5), .ZN(n946) );
  NAND2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G21), .B(G1966), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(KEYINPUT127), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(KEYINPUT61), .B(n953), .Z(n954) );
  NOR2_X1 U1054 ( .A1(G16), .A2(n954), .ZN(n982) );
  XNOR2_X1 U1055 ( .A(KEYINPUT56), .B(G16), .ZN(n979) );
  XNOR2_X1 U1056 ( .A(n956), .B(n955), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(KEYINPUT57), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G301), .B(G1961), .ZN(n964) );
  XOR2_X1 U1062 ( .A(n962), .B(G1348), .Z(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1064 ( .A(KEYINPUT122), .B(n965), .Z(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G1956), .B(G299), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(KEYINPUT123), .B(n980), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n1013) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT120), .B(n983), .ZN(n986) );
  XOR2_X1 U1078 ( .A(G2072), .B(n984), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT50), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n996) );
  XOR2_X1 U1082 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n994) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT118), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1007) );
  XNOR2_X1 U1088 ( .A(G160), .B(G2084), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT117), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT121), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1009), .ZN(n1010) );
  INV_X1 U1097 ( .A(KEYINPUT55), .ZN(n1032) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1032), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(G29), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1037) );
  XNOR2_X1 U1101 ( .A(G2090), .B(G35), .ZN(n1027) );
  XNOR2_X1 U1102 ( .A(G1996), .B(G32), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G33), .B(G2072), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(G25), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(G28), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G26), .B(G2067), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(G27), .B(n1022), .Z(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT53), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(G2084), .B(G34), .Z(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT54), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(n1032), .B(n1031), .ZN(n1034) );
  INV_X1 U1118 ( .A(G29), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(G11), .A2(n1035), .ZN(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(n1038), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

