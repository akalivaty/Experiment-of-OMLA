//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n643, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n464), .B2(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(KEYINPUT68), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n479), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n464), .A2(new_n465), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(G114), .B2(new_n463), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n464), .B2(new_n465), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n505), .C1(new_n465), .C2(new_n464), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n475), .A2(new_n479), .A3(new_n508), .A4(new_n502), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n500), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT73), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(KEYINPUT72), .A3(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n516), .A2(KEYINPUT74), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT74), .B1(new_n516), .B2(new_n525), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NOR3_X1   g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI211_X1 g104(.A(new_n511), .B(new_n521), .C1(new_n523), .C2(new_n524), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT75), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n513), .B1(new_n514), .B2(G543), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n511), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n521), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n520), .A2(KEYINPUT72), .A3(G651), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT72), .B1(new_n520), .B2(G651), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n534), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n516), .A2(new_n525), .A3(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G88), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(new_n546), .A3(new_n531), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n519), .B1(new_n533), .B2(new_n547), .ZN(G166));
  NOR2_X1   g123(.A1(new_n526), .A2(new_n527), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n530), .A2(G51), .B1(new_n516), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n549), .A2(G89), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT7), .Z(new_n555));
  NAND2_X1  g130(.A1(new_n516), .A2(new_n550), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n525), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G51), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n555), .B1(new_n559), .B2(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n553), .A2(new_n560), .ZN(G286));
  INV_X1    g136(.A(G286), .ZN(G168));
  AND2_X1   g137(.A1(G77), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n516), .B2(G64), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n518), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  XNOR2_X1  g141(.A(KEYINPUT78), .B(G52), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n566), .B1(new_n530), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT79), .B(G90), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n549), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n564), .B2(new_n518), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(G301));
  INV_X1    g147(.A(G301), .ZN(G171));
  NAND2_X1  g148(.A1(new_n549), .A2(G81), .ZN(new_n574));
  NAND2_X1  g149(.A1(G68), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G56), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n538), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G43), .B2(new_n530), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G860), .ZN(G153));
  NAND4_X1  g156(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT8), .ZN(new_n585));
  NAND4_X1  g160(.A1(G319), .A2(G483), .A3(G661), .A4(new_n585), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT81), .Z(G188));
  NAND2_X1  g162(.A1(new_n523), .A2(new_n524), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n588), .A2(G53), .A3(G543), .A4(new_n539), .ZN(new_n589));
  NAND2_X1  g164(.A1(KEYINPUT82), .A2(KEYINPUT9), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n525), .A2(G53), .A3(G543), .A4(new_n590), .ZN(new_n593));
  OAI211_X1 g168(.A(G65), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n594));
  NAND2_X1  g169(.A1(G78), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n592), .A2(new_n593), .B1(new_n596), .B2(G651), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n543), .A2(G91), .A3(new_n544), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G299));
  INV_X1    g174(.A(new_n519), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n545), .A2(new_n546), .A3(new_n531), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n546), .B1(new_n545), .B2(new_n531), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(G303));
  OR2_X1    g178(.A1(new_n516), .A2(G74), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G49), .B2(new_n530), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n543), .A2(G87), .A3(new_n544), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G288));
  NAND2_X1  g182(.A1(G73), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n538), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G48), .B2(new_n530), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n543), .A2(G86), .A3(new_n544), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G305));
  AOI22_X1  g188(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n518), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n530), .A2(G47), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n543), .A2(new_n544), .ZN(new_n617));
  INV_X1    g192(.A(G85), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g196(.A(KEYINPUT83), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n549), .A2(KEYINPUT10), .A3(G92), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(G79), .A2(G543), .ZN(new_n631));
  INV_X1    g206(.A(G66), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n538), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n633), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n625), .B1(new_n636), .B2(G868), .ZN(G284));
  XOR2_X1   g212(.A(G284), .B(KEYINPUT84), .Z(G321));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(G299), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G168), .B2(new_n639), .ZN(G297));
  OAI21_X1  g216(.A(new_n640), .B1(G168), .B2(new_n639), .ZN(G280));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n636), .B1(new_n643), .B2(G860), .ZN(G148));
  NOR2_X1   g219(.A1(new_n579), .A2(G868), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n636), .A2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n645), .B1(new_n647), .B2(G868), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n487), .A2(G123), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n463), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(G135), .B2(new_n485), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n475), .A2(new_n479), .A3(new_n469), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G2100), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(G2100), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(G156));
  XOR2_X1   g238(.A(KEYINPUT15), .B(G2435), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(KEYINPUT14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2451), .B(G2454), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n678), .A2(new_n679), .A3(G14), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT89), .ZN(G401));
  XOR2_X1   g256(.A(G2067), .B(G2678), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT18), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n684), .B(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n686), .C1(new_n683), .C2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n683), .A3(new_n685), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2096), .B(G2100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1971), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n698), .B2(new_n704), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT92), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(G229));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G1966), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(G1966), .ZN(new_n720));
  NOR2_X1   g295(.A1(G4), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n636), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1348), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n655), .A2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT103), .ZN(new_n726));
  NOR2_X1   g301(.A1(G29), .A2(G35), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G162), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G28), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT30), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n732), .B2(KEYINPUT30), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  INV_X1    g314(.A(G129), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n498), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n485), .A2(G141), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n469), .A2(G105), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n746), .B2(G32), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT27), .B(G1996), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT101), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n737), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n750), .B2(new_n748), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n726), .A2(new_n731), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n580), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G19), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT96), .B(G1341), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n746), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n485), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n487), .A2(G128), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n765), .A2(KEYINPUT97), .A3(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT97), .B1(new_n765), .B2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n757), .A2(new_n758), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n746), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n746), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(G29), .A2(G33), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n485), .A2(G139), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT98), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n475), .A2(new_n479), .A3(G127), .ZN(new_n781));
  NAND2_X1  g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n778), .B(new_n780), .C1(new_n783), .C2(new_n463), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(new_n746), .ZN(new_n785));
  INV_X1    g360(.A(G2072), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n785), .A2(new_n786), .B1(new_n774), .B2(new_n773), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n775), .B(new_n787), .C1(new_n786), .C2(new_n785), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n753), .A2(new_n771), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G34), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(KEYINPUT24), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(KEYINPUT24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n746), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G160), .B2(new_n746), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT99), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2084), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT104), .B(KEYINPUT23), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT105), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n715), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  INV_X1    g376(.A(G299), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n715), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n797), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n715), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n715), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1961), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  INV_X1    g384(.A(new_n795), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n724), .A2(new_n789), .A3(new_n805), .A4(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT106), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n715), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n623), .B2(new_n715), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n485), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n487), .A2(G119), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n463), .A2(G107), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT93), .Z(new_n823));
  MUX2_X1   g398(.A(G25), .B(new_n823), .S(G29), .Z(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G288), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n715), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n715), .B2(G23), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT95), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G22), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G166), .B2(G16), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n833), .B(new_n837), .C1(G1971), .C2(new_n839), .ZN(new_n840));
  MUX2_X1   g415(.A(G6), .B(G305), .S(G16), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT94), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT32), .B(G1981), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G1971), .ZN(new_n845));
  INV_X1    g420(.A(new_n839), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT34), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n827), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT34), .B1(new_n840), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT36), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT36), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n814), .B1(new_n853), .B2(new_n855), .ZN(G311));
  XNOR2_X1  g431(.A(new_n812), .B(KEYINPUT106), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n854), .B1(new_n850), .B2(new_n851), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G150));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n617), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G55), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n863), .A2(new_n518), .B1(new_n864), .B2(new_n557), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT110), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT108), .B1(new_n579), .B2(KEYINPUT107), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n574), .A2(new_n872), .A3(new_n873), .A4(new_n578), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n867), .B1(new_n580), .B2(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n866), .B1(new_n579), .B2(KEYINPUT107), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n871), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n635), .A2(new_n643), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT39), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT109), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT39), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(G860), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n870), .B1(new_n887), .B2(new_n889), .ZN(G145));
  XNOR2_X1  g465(.A(new_n784), .B(new_n745), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n487), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n463), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G142), .B2(new_n485), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(new_n658), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n891), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G164), .B(new_n765), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n822), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(G160), .B(G162), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n655), .ZN(new_n903));
  AOI21_X1  g478(.A(G37), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n903), .B2(new_n901), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g481(.A1(new_n647), .A2(new_n879), .A3(new_n877), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT85), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n646), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n880), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n635), .A2(G299), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n630), .A2(new_n802), .A3(new_n634), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n907), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n907), .A2(new_n910), .ZN(new_n920));
  INV_X1    g495(.A(new_n913), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n907), .A2(new_n910), .A3(new_n917), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n907), .B2(new_n910), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n623), .A2(G303), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G288), .B(G305), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n623), .A2(G303), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n934), .A2(KEYINPUT111), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n922), .A2(new_n925), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n922), .B2(new_n925), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n867), .A2(new_n639), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  XOR2_X1   g516(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  AND2_X1   g519(.A1(G286), .A2(G301), .ZN(new_n945));
  NOR2_X1   g520(.A1(G286), .A2(G301), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n877), .A2(new_n947), .A3(new_n879), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n879), .B2(new_n877), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n949), .A3(new_n913), .ZN(new_n950));
  INV_X1    g525(.A(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n880), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n877), .A2(new_n947), .A3(new_n879), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n917), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n944), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n921), .A3(new_n953), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n948), .A2(new_n949), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(KEYINPUT113), .C1(new_n957), .C2(new_n917), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n934), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n933), .B(new_n956), .C1(new_n957), .C2(new_n917), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n943), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n934), .B1(new_n950), .B2(new_n954), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n961), .A3(new_n960), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n942), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n965), .A2(new_n968), .A3(KEYINPUT43), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(new_n962), .A3(new_n943), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n971), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT127), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n765), .A2(G2067), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n505), .B1(new_n497), .B2(new_n502), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n509), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G114), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n494), .B1(new_n980), .B2(G2105), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n487), .B2(G126), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT115), .B(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n480), .A2(new_n481), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G2105), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n466), .A2(new_n470), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT69), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n993), .A3(G40), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n765), .B(G2067), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n745), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n745), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(G1996), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n825), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n823), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n976), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n996), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT125), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n822), .B(new_n1007), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n995), .A2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1006), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(G290), .A2(new_n996), .A3(G1986), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT48), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n995), .B1(new_n1001), .B2(new_n997), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n996), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n995), .B2(new_n998), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1012), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n975), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1027), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(KEYINPUT127), .A3(new_n1012), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n983), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n994), .B1(new_n1035), .B2(new_n986), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n983), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n983), .A2(new_n1040), .A3(new_n1034), .ZN(new_n1041));
  INV_X1    g616(.A(G40), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n473), .A2(new_n482), .A3(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(new_n809), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1033), .B1(new_n1046), .B2(KEYINPUT122), .ZN(new_n1047));
  OAI21_X1  g622(.A(G286), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n986), .B1(G164), .B2(G1384), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1050));
  INV_X1    g625(.A(G1966), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(G168), .A3(new_n1044), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1053), .A3(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1052), .B2(new_n1044), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT51), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1053), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n983), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1049), .A2(new_n1063), .A3(new_n1043), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1049), .A2(new_n1063), .A3(new_n1066), .A4(new_n1043), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n845), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n994), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(new_n730), .A3(new_n1041), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1056), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(G166), .A2(new_n1056), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(G303), .B2(G8), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n611), .A2(new_n1079), .A3(new_n612), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n611), .B2(new_n612), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n611), .A2(new_n1079), .A3(new_n612), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT49), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G164), .A2(G1384), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1056), .B1(new_n1086), .B2(new_n1043), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n605), .A2(new_n606), .A3(G1976), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT52), .ZN(new_n1091));
  INV_X1    g666(.A(G1976), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1088), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1062), .A2(new_n1077), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n597), .A2(new_n1099), .A3(new_n598), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n597), .B2(new_n598), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1049), .A2(new_n1063), .A3(new_n1043), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1035), .A2(new_n994), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1103), .A2(new_n1109), .B1(new_n1110), .B2(new_n769), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n635), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT61), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1102), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1956), .B1(new_n1069), .B2(new_n1041), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1107), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1113), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1113), .A3(new_n1115), .A4(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1111), .A2(new_n1124), .A3(new_n636), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1110), .A2(new_n769), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1126), .A2(new_n635), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1049), .A2(new_n1063), .A3(new_n998), .A4(new_n1043), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1035), .B2(new_n994), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1132), .B1(new_n1136), .B2(new_n580), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1132), .A3(new_n580), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1131), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT120), .B(new_n579), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1137), .A2(new_n1141), .A3(KEYINPUT59), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1114), .B1(new_n1130), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n774), .A2(KEYINPUT53), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n987), .A2(new_n1043), .A3(new_n1063), .A4(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g722(.A(G1961), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1103), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(G2078), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1147), .B(new_n1149), .C1(KEYINPUT53), .C2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G301), .B(KEYINPUT54), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1036), .A2(new_n1037), .A3(new_n1145), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n1149), .C1(new_n1150), .C2(KEYINPUT53), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1156), .B2(new_n1153), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1098), .A2(new_n1144), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1077), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n1096), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1055), .A2(new_n1161), .A3(new_n1061), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1156), .A2(G171), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1159), .A2(new_n1096), .A3(new_n1164), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1169), .B2(new_n1162), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1158), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(G8), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1046), .A2(G286), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1077), .A3(new_n1095), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1097), .A2(KEYINPUT63), .A3(new_n1077), .A4(new_n1176), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1088), .A2(new_n1092), .A3(new_n828), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1087), .B1(new_n1182), .B2(new_n1080), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1095), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT119), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1188), .B(new_n1185), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1171), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n623), .B(G1986), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1015), .B1(new_n996), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1032), .B1(new_n1190), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(new_n461), .ZN(new_n1195));
  NOR4_X1   g769(.A1(G229), .A2(new_n1195), .A3(new_n680), .A4(G227), .ZN(new_n1196));
  OAI211_X1 g770(.A(new_n1196), .B(new_n905), .C1(new_n963), .C2(new_n966), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


