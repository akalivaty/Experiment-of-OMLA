//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n205), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AND2_X1   g0018(.A1(KEYINPUT64), .A2(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(KEYINPUT64), .A2(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n213), .A2(new_n216), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n212), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT67), .Z(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G222), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n249), .B1(new_n250), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n259), .A2(G274), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT68), .A2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT68), .A2(G45), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n255), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n256), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g0075(.A(KEYINPUT8), .B(G58), .Z(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G33), .A3(new_n221), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n202), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  INV_X1    g0084(.A(G20), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n284), .A2(new_n285), .A3(G1), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n240), .B1(new_n265), .B2(G20), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n287), .A2(new_n288), .B1(new_n240), .B2(new_n286), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n256), .A2(new_n268), .A3(new_n272), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n275), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n265), .A2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n287), .A2(G77), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n284), .A2(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G20), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(G77), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n281), .A2(new_n222), .ZN(new_n302));
  OR2_X1    g0102(.A1(KEYINPUT64), .A2(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT64), .A2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n276), .A2(new_n278), .B1(new_n305), .B2(G77), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G33), .A3(new_n221), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n248), .A2(G232), .A3(new_n251), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G107), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n248), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n255), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n271), .A2(G244), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n268), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n311), .B1(new_n318), .B2(new_n292), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G179), .B2(new_n318), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n311), .C1(new_n322), .C2(new_n318), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n296), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n290), .B(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n273), .A2(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n291), .A2(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT10), .Z(new_n329));
  INV_X1    g0129(.A(KEYINPUT72), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n248), .A2(G232), .A3(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n332), .A2(new_n334), .A3(G226), .A4(new_n251), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n255), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n271), .A2(G238), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n268), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n342));
  NAND4_X1  g0142(.A1(new_n268), .A2(new_n338), .A3(new_n342), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(G190), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n242), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n221), .A2(G33), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n250), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n282), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT11), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n300), .A2(KEYINPUT12), .A3(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT12), .B1(new_n300), .B2(G68), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n242), .B1(new_n265), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n352), .A2(new_n353), .B1(new_n287), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  INV_X1    g0159(.A(new_n342), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n340), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n330), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n262), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT68), .A2(G45), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n364), .A2(new_n365), .A3(G41), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT69), .B1(new_n366), .B2(G1), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n260), .B1(G238), .B2(new_n271), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n342), .B1(new_n370), .B2(new_n338), .ZN(new_n371));
  INV_X1    g0171(.A(new_n343), .ZN(new_n372));
  OAI21_X1  g0172(.A(G200), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT72), .A3(new_n344), .A4(new_n357), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(G169), .C1(new_n371), .C2(new_n372), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n341), .A2(G179), .A3(new_n343), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n361), .A2(new_n343), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(G169), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n356), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n324), .A2(new_n329), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n287), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n276), .A2(new_n297), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n385), .A2(new_n386), .B1(new_n300), .B2(new_n276), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT75), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n332), .A2(new_n334), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n285), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT74), .ZN(new_n394));
  AOI21_X1  g0194(.A(G20), .B1(new_n332), .B2(new_n334), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT7), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT73), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT73), .B1(new_n332), .B2(new_n334), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n398), .A2(new_n399), .A3(new_n305), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n394), .B(new_n397), .C1(new_n400), .C2(KEYINPUT7), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n391), .B1(new_n401), .B2(G68), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n302), .B1(new_n402), .B2(KEYINPUT16), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT7), .B1(new_n305), .B2(new_n248), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n390), .B1(new_n407), .B2(new_n242), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n388), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G87), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n257), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n392), .A2(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(G223), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n332), .A2(new_n334), .A3(G226), .A4(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT76), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n248), .A2(new_n418), .A3(G226), .A4(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n255), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n271), .A2(G232), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(G179), .A3(new_n268), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n268), .A2(new_n423), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n259), .B1(new_n415), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT18), .B1(new_n411), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n398), .A2(new_n399), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT7), .B1(new_n431), .B2(new_n221), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n394), .A2(new_n397), .ZN(new_n433));
  OAI21_X1  g0233(.A(G68), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT16), .A3(new_n390), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n410), .A3(new_n282), .ZN(new_n436));
  INV_X1    g0236(.A(new_n388), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n428), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n359), .B1(new_n425), .B2(new_n426), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n422), .A2(new_n268), .A3(new_n423), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(G190), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n436), .A2(new_n444), .A3(new_n437), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n436), .A2(new_n444), .A3(KEYINPUT17), .A4(new_n437), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(KEYINPUT77), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n430), .A2(new_n440), .A3(new_n447), .A4(new_n448), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n384), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n332), .A2(new_n334), .A3(G257), .A4(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n332), .A2(new_n334), .A3(G250), .A4(new_n251), .ZN(new_n457));
  INV_X1    g0257(.A(G294), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n257), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n265), .A2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n258), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n255), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n459), .A2(new_n255), .B1(new_n465), .B2(G264), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(G274), .A3(new_n259), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n292), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G179), .B2(new_n468), .ZN(new_n470));
  XOR2_X1   g0270(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n221), .A2(new_n248), .A3(G87), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n474), .A2(G87), .A3(new_n221), .A4(new_n248), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n314), .C1(new_n219), .C2(new_n220), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n479), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n285), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT23), .A2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n472), .B1(new_n478), .B2(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n471), .B(new_n485), .C1(new_n476), .C2(new_n477), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n282), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT88), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT88), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n282), .C1(new_n487), .C2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n314), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT25), .B1(new_n286), .B2(new_n314), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n265), .A2(G33), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n302), .A2(new_n300), .A3(new_n497), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n495), .A2(new_n496), .B1(new_n498), .B2(new_n314), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n470), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n459), .A2(new_n255), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n465), .A2(G264), .ZN(new_n503));
  AND4_X1   g0303(.A1(new_n322), .A2(new_n502), .A3(new_n503), .A4(new_n467), .ZN(new_n504));
  AOI21_X1  g0304(.A(G200), .B1(new_n466), .B2(new_n467), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n499), .B(new_n506), .C1(new_n490), .C2(new_n492), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT89), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n506), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n493), .A2(new_n500), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT89), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n499), .B1(new_n490), .B2(new_n492), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n511), .C1(new_n512), .C2(new_n470), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT79), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  INV_X1    g0316(.A(new_n278), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n250), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n278), .A2(KEYINPUT78), .A3(G77), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g0320(.A(G97), .B(G107), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n522), .A2(new_n524), .A3(G107), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n520), .B1(new_n527), .B2(new_n305), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n404), .A2(new_n406), .A3(G107), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n302), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n300), .A2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n498), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n515), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n529), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n525), .B1(new_n522), .B2(new_n521), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n518), .B(new_n519), .C1(new_n537), .C2(new_n221), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n282), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(KEYINPUT79), .A3(new_n533), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n465), .A2(new_n542), .A3(G257), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n269), .A2(G1), .ZN(new_n544));
  INV_X1    g0344(.A(new_n463), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(G257), .A3(new_n259), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n543), .A2(new_n549), .B1(new_n260), .B2(new_n464), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n332), .A2(new_n334), .A3(G244), .A4(new_n251), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n332), .A2(new_n334), .A3(G250), .A4(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n551), .C2(new_n552), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT80), .B1(new_n551), .B2(new_n552), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n550), .B(new_n322), .C1(new_n259), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n543), .A2(new_n549), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n467), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n259), .B1(new_n563), .B2(new_n553), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n560), .B1(new_n565), .B2(G200), .ZN(new_n566));
  OAI21_X1  g0366(.A(G169), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n550), .B(G179), .C1(new_n259), .C2(new_n559), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n539), .A2(new_n533), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n541), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n303), .A2(new_n304), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT82), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n221), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n412), .A2(new_n524), .A3(new_n314), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n303), .A2(G33), .A3(G97), .A4(new_n304), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n221), .A2(new_n248), .A3(G68), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n282), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n498), .A2(new_n307), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n308), .A2(new_n300), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n582), .A3(new_n581), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n593), .B2(new_n282), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(KEYINPUT83), .A3(new_n586), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n460), .A2(G250), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n260), .A2(new_n544), .B1(new_n259), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n332), .A2(new_n334), .A3(G238), .A4(new_n251), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n332), .A2(new_n334), .A3(G244), .A4(G1698), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n481), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n255), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(G179), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n292), .B2(new_n603), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n602), .A3(G190), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n532), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n603), .A2(G200), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n594), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n596), .A2(new_n605), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n257), .A2(G97), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n303), .A2(new_n613), .A3(new_n304), .A4(new_n556), .ZN(new_n614));
  INV_X1    g0414(.A(G116), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n281), .A2(new_n222), .B1(G20), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n498), .B2(new_n615), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n287), .A2(KEYINPUT85), .A3(G116), .A4(new_n497), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n286), .A2(new_n615), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n547), .A2(G270), .A3(new_n259), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n467), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n332), .A2(new_n334), .A3(G264), .A4(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n332), .A2(new_n334), .A3(G257), .A4(new_n251), .ZN(new_n629));
  INV_X1    g0429(.A(G303), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n248), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n255), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n292), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n619), .A2(new_n624), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n627), .A2(new_n632), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G200), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n627), .A2(new_n632), .A3(G190), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n623), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n467), .A2(new_n626), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n255), .B2(new_n631), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n625), .A2(G179), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n625), .A2(KEYINPUT21), .A3(new_n633), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n636), .A2(new_n641), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n571), .A2(new_n612), .A3(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n455), .A2(new_n514), .A3(new_n647), .ZN(G372));
  INV_X1    g0448(.A(KEYINPUT90), .ZN(new_n649));
  INV_X1    g0449(.A(new_n382), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n320), .B1(new_n363), .B2(new_n374), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n449), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n650), .A2(new_n651), .A3(new_n649), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n441), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n328), .A2(KEYINPUT10), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n328), .A2(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n296), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n571), .A2(new_n510), .A3(new_n612), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n636), .A2(new_n644), .A3(new_n645), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n493), .A2(new_n500), .ZN(new_n663));
  INV_X1    g0463(.A(new_n470), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT83), .B1(new_n594), .B2(new_n586), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n581), .A2(new_n582), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n302), .B1(new_n668), .B2(new_n592), .ZN(new_n669));
  NOR4_X1   g0469(.A1(new_n669), .A2(new_n590), .A3(new_n585), .A4(new_n587), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n605), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n611), .A2(new_n608), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n569), .A2(new_n570), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n567), .A2(new_n568), .B1(new_n535), .B2(new_n540), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n671), .A3(new_n677), .A4(new_n672), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n671), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n666), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n454), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n660), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n221), .A2(new_n299), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  INV_X1    g0485(.A(G213), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n683), .B2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n514), .B1(new_n663), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n501), .B2(new_n690), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n690), .A2(new_n625), .ZN(new_n693));
  MUX2_X1   g0493(.A(new_n646), .B(new_n662), .S(new_n693), .Z(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n662), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n514), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n512), .A2(new_n470), .A3(new_n690), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0507(.A(new_n214), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n577), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n218), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n680), .A2(new_n701), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n535), .A2(new_n540), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n569), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT26), .B1(new_n673), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n569), .A2(new_n570), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n612), .A2(new_n677), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n723), .A3(new_n671), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n701), .C1(new_n666), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n597), .A2(new_n259), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n259), .A2(G274), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n460), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n255), .B2(new_n601), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n643), .A2(new_n732), .A3(G179), .A4(new_n466), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n550), .B1(new_n559), .B2(new_n259), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n728), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n502), .A2(new_n598), .A3(new_n602), .A4(new_n503), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n627), .A2(new_n632), .A3(G179), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n728), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n565), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n732), .A2(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n734), .A2(new_n468), .A3(new_n741), .A4(new_n638), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n735), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n690), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n571), .A2(new_n612), .A3(new_n646), .A4(new_n701), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n747), .C1(new_n514), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n726), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n715), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n305), .A2(new_n284), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G45), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G1), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n709), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n695), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n322), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n221), .B1(new_n274), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n392), .B1(new_n764), .B2(new_n458), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n359), .A2(G179), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n285), .A2(new_n322), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n221), .A2(new_n274), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n322), .A3(new_n359), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n630), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n763), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n765), .B(new_n773), .C1(G322), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n770), .A2(G200), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n778), .B2(new_n322), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(KEYINPUT96), .A3(G190), .A4(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n778), .A2(G190), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n784));
  INV_X1    g0584(.A(G317), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n221), .A2(KEYINPUT97), .A3(G190), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT97), .B1(new_n221), .B2(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(new_n767), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G283), .A2(new_n791), .B1(new_n794), .B2(G329), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n776), .A2(new_n782), .A3(new_n787), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n769), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G87), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n775), .A2(G58), .ZN(new_n799));
  INV_X1    g0599(.A(new_n764), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G97), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n798), .A2(new_n799), .A3(new_n248), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G68), .B2(new_n783), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G77), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n781), .A2(G50), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n791), .A2(G107), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n803), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n794), .A2(G159), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT32), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n796), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n222), .B1(G20), .B2(new_n292), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n761), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n431), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n708), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n261), .A2(new_n262), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n713), .B2(new_n819), .C1(new_n246), .C2(new_n269), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n708), .A2(new_n392), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G355), .B1(new_n615), .B2(new_n708), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n758), .B1(new_n762), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n694), .B(G330), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n758), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT100), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  OAI21_X1  g0629(.A(new_n323), .B1(new_n701), .B2(new_n311), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n320), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n320), .A2(new_n690), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n716), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n701), .B(new_n835), .C1(new_n666), .C2(new_n679), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n757), .B1(new_n837), .B2(new_n750), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n750), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n815), .A2(new_n759), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n758), .B1(new_n250), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n791), .A2(G87), .ZN(new_n842));
  INV_X1    g0642(.A(new_n783), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n846), .A2(G283), .B1(G303), .B2(new_n781), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n801), .B(new_n392), .C1(new_n314), .C2(new_n769), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G294), .B2(new_n775), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n807), .A2(G116), .B1(G311), .B2(new_n794), .ZN(new_n850));
  AND4_X1   g0650(.A1(new_n842), .A2(new_n847), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n843), .A2(new_n852), .B1(new_n853), .B2(new_n774), .ZN(new_n854));
  INV_X1    g0654(.A(G159), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n806), .A2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G137), .C2(new_n781), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n791), .A2(G68), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n794), .A2(G132), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n797), .A2(G50), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n431), .B1(new_n800), .B2(G58), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n815), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n841), .B1(new_n760), .B2(new_n835), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n839), .A2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n754), .A2(new_n265), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  INV_X1    g0671(.A(new_n688), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT37), .B1(new_n438), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n438), .A2(new_n428), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n445), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n248), .A2(KEYINPUT74), .A3(new_n405), .A4(G20), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n396), .B1(new_n395), .B2(KEYINPUT7), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT73), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n392), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT73), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n221), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n405), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n242), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n409), .B1(new_n885), .B2(new_n391), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n387), .B1(new_n403), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n424), .A2(new_n427), .A3(new_n688), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n445), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT37), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n876), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n435), .A3(new_n282), .ZN(new_n896));
  INV_X1    g0696(.A(new_n387), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n451), .A2(new_n872), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n871), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n888), .ZN(new_n902));
  AOI211_X1 g0702(.A(KEYINPUT102), .B(new_n901), .C1(new_n902), .C2(new_n445), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n893), .B1(new_n890), .B2(KEYINPUT37), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n875), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n451), .A2(new_n872), .A3(new_n898), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n690), .A2(new_n356), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n375), .A2(new_n382), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n375), .B2(new_n382), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n835), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n508), .A2(new_n513), .ZN(new_n914));
  INV_X1    g0714(.A(new_n748), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n746), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n912), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT40), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT104), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n445), .B1(new_n411), .B2(new_n429), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n901), .B1(new_n411), .B2(new_n688), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n873), .A2(KEYINPUT104), .A3(new_n874), .A4(new_n445), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n411), .A2(new_n688), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT37), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n451), .A2(new_n438), .A3(new_n872), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n907), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n748), .B1(new_n508), .B2(new_n513), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n936), .A2(new_n919), .A3(new_n913), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n912), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n922), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n455), .A2(new_n937), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n696), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n945));
  INV_X1    g0745(.A(new_n933), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n930), .B2(new_n931), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n650), .A2(new_n701), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n441), .A2(new_n872), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n910), .A2(new_n911), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n836), .B2(new_n832), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n953), .B1(new_n908), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n718), .A2(new_n454), .A3(new_n725), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n660), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n870), .B1(new_n943), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n943), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n963), .A2(G116), .A3(new_n223), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  INV_X1    g0766(.A(G58), .ZN(new_n967));
  OAI21_X1  g0767(.A(G77), .B1(new_n967), .B2(new_n242), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n241), .B1(new_n713), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n284), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n966), .A3(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n571), .B1(new_n541), .B2(new_n701), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n676), .A2(new_n690), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT106), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n699), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n501), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n701), .B1(new_n977), .B2(new_n722), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n703), .A2(new_n974), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(KEYINPUT107), .A3(new_n980), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(KEYINPUT42), .C2(new_n979), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n594), .A2(new_n609), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n612), .B1(new_n986), .B2(new_n701), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n671), .A2(new_n986), .A3(new_n701), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n985), .B2(new_n992), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n976), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n995), .ZN(new_n997));
  INV_X1    g0797(.A(new_n976), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(new_n993), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n709), .B(KEYINPUT41), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n705), .A2(new_n974), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n705), .A2(new_n974), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n700), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n699), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n692), .A2(new_n702), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n514), .B2(new_n702), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n697), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n698), .C1(new_n514), .C2(new_n702), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n751), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1009), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1000), .B1(new_n1017), .B2(new_n752), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n996), .B(new_n999), .C1(new_n756), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n761), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n989), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n846), .A2(G159), .B1(G143), .B2(new_n781), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n790), .A2(new_n250), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n800), .A2(G68), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n248), .C1(new_n967), .C2(new_n769), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(G150), .C2(new_n775), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n807), .A2(G50), .B1(G137), .B2(new_n794), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n431), .B1(new_n764), .B2(new_n314), .C1(new_n774), .C2(new_n630), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n806), .A2(new_n1030), .B1(new_n785), .B2(new_n793), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G97), .C2(new_n791), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n769), .A2(new_n615), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT46), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n846), .B2(G294), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n781), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1032), .B1(KEYINPUT109), .B2(new_n1035), .C1(new_n772), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(KEYINPUT109), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1028), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT47), .Z(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n867), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n818), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n816), .B1(new_n214), .B2(new_n307), .C1(new_n1042), .C2(new_n235), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT108), .Z(new_n1044));
  NOR3_X1   g0844(.A1(new_n1041), .A2(new_n758), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT110), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1021), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1019), .A2(new_n1048), .ZN(G387));
  OAI22_X1  g0849(.A1(new_n769), .A2(new_n250), .B1(new_n774), .B2(new_n240), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n800), .A2(new_n308), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n817), .C1(new_n242), .C2(new_n771), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n276), .C2(new_n783), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G97), .A2(new_n791), .B1(new_n794), .B2(G150), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n781), .A2(KEYINPUT111), .A3(G159), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT111), .B1(new_n781), .B2(G159), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1054), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n817), .B1(new_n794), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n769), .A2(new_n458), .B1(new_n1030), .B2(new_n764), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n807), .A2(G303), .B1(G317), .B2(new_n775), .ZN(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n846), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1036), .C1(new_n1062), .C2(new_n772), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1058), .B1(new_n615), .B2(new_n790), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1057), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n815), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n231), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1042), .B1(new_n1072), .B2(new_n819), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n711), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n821), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n711), .B(new_n269), .C1(new_n242), .C2(new_n250), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n276), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(G50), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n276), .A2(KEYINPUT50), .A3(new_n240), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1075), .A2(new_n1081), .B1(G107), .B2(new_n214), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n758), .B1(new_n1082), .B2(new_n816), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1071), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n692), .B2(new_n761), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n756), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1016), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n709), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1086), .A2(new_n752), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  AOI21_X1  g0891(.A(new_n700), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1010), .A2(new_n699), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n756), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n816), .B1(new_n524), .B2(new_n214), .C1(new_n1042), .C2(new_n239), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1096), .A2(new_n757), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n793), .A2(new_n1061), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n771), .A2(new_n458), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n797), .A2(G283), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n248), .B1(new_n800), .B2(G116), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n810), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(G303), .C2(new_n846), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n781), .A2(G317), .B1(G311), .B2(new_n775), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n797), .A2(G68), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n800), .A2(G77), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n842), .A2(new_n817), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n806), .A2(new_n1078), .B1(new_n853), .B2(new_n793), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G50), .C2(new_n846), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n781), .A2(G150), .B1(G159), .B2(new_n775), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT51), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1106), .B1(new_n1115), .B2(KEYINPUT112), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT112), .B2(new_n1115), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1097), .B1(new_n975), .B2(new_n1020), .C1(new_n867), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1094), .A2(new_n1016), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1017), .A2(new_n709), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1095), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n916), .A2(new_n920), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n454), .A2(G330), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n660), .A2(new_n958), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n912), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(G330), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT113), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n749), .A2(G330), .A3(new_n835), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n954), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1122), .A2(KEYINPUT113), .A3(new_n1125), .A4(G330), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n836), .A2(new_n832), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n701), .B(new_n831), .C1(new_n666), .C2(new_n724), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n832), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1129), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n954), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1122), .A2(G330), .A3(new_n835), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n954), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1124), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n950), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n948), .B2(new_n951), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n935), .A2(new_n1148), .A3(new_n949), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n949), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT38), .B1(new_n905), .B2(new_n906), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n945), .A2(new_n1153), .A3(new_n944), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT39), .B1(new_n934), .B2(new_n907), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n935), .A2(new_n1148), .A3(new_n949), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1150), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1144), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1124), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n1159), .A3(new_n1150), .A4(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n709), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n756), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n759), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n840), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n757), .B1(new_n276), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n846), .A2(G107), .B1(G283), .B2(new_n781), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n798), .A2(new_n392), .A3(new_n1108), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G116), .B2(new_n775), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n807), .A2(G97), .B1(G294), .B2(new_n794), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n859), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT114), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT114), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n797), .A2(G150), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT54), .B(G143), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n807), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n240), .B2(new_n790), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n392), .B1(new_n800), .B2(G159), .ZN(new_n1183));
  INV_X1    g0983(.A(G132), .ZN(new_n1184));
  INV_X1    g0984(.A(G125), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1183), .B1(new_n774), .B2(new_n1184), .C1(new_n793), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n781), .B2(G128), .ZN(new_n1187));
  INV_X1    g0987(.A(G137), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1062), .B2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1176), .B(new_n1177), .C1(new_n1182), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1170), .B1(new_n1190), .B2(new_n815), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1167), .B1(new_n1168), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n1192), .ZN(G378));
  NOR2_X1   g0993(.A1(new_n945), .A2(new_n947), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1122), .A2(KEYINPUT40), .A3(new_n1125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(G330), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n688), .B1(new_n283), .B2(new_n289), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n294), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n329), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1197), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n658), .A2(new_n294), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1200), .B1(new_n658), .B2(new_n294), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1198), .B(new_n1197), .C1(new_n656), .C2(new_n657), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT116), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n1207), .A3(KEYINPUT116), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1196), .A2(new_n922), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n921), .B1(new_n945), .B2(new_n1153), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n938), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n696), .B1(new_n939), .B2(new_n935), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n957), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n957), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1208), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1196), .B2(new_n922), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1212), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n756), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n757), .B1(G50), .B2(new_n1169), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1024), .B1(new_n250), .B2(new_n769), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n817), .A2(G41), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n314), .B2(new_n774), .C1(new_n307), .C2(new_n771), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G97), .C2(new_n783), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n790), .A2(new_n967), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G283), .B2(new_n794), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(new_n615), .C2(new_n1036), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT58), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1229), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G50), .B1(new_n257), .B2(new_n258), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1234), .A2(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n797), .A2(new_n1180), .B1(new_n775), .B2(G128), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT115), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n771), .A2(new_n1188), .B1(new_n852), .B2(new_n764), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G132), .B2(new_n783), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n1185), .C2(new_n1036), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n257), .B(new_n258), .C1(new_n790), .C2(new_n855), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G124), .B2(new_n794), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1238), .B1(new_n1235), .B2(new_n1234), .C1(new_n1244), .C2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1227), .B1(new_n1249), .B2(new_n815), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1222), .B2(new_n760), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1164), .A2(new_n1163), .B1(new_n1224), .B2(new_n1218), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n709), .B1(new_n1253), .B2(KEYINPUT57), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT117), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1218), .A2(new_n1224), .A3(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1133), .A2(new_n1132), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1163), .B1(new_n1160), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1219), .A2(new_n1223), .A3(new_n1221), .A4(KEYINPUT117), .ZN(new_n1259));
  AND4_X1   g1059(.A1(KEYINPUT57), .A2(new_n1256), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1254), .B2(new_n1260), .ZN(G375));
  INV_X1    g1061(.A(new_n1000), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1134), .A2(new_n1142), .A3(new_n1124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1144), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n954), .A2(new_n759), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT118), .Z(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n757), .B1(G68), .B2(new_n1169), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n846), .A2(new_n1180), .B1(G137), .B2(new_n775), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1184), .B2(new_n1036), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT120), .Z(new_n1271));
  AOI21_X1  g1071(.A(new_n431), .B1(new_n800), .B2(G50), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n852), .B2(new_n771), .C1(new_n855), .C2(new_n769), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n794), .A2(G128), .ZN(new_n1274));
  OR3_X1    g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1232), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n793), .A2(new_n630), .B1(new_n769), .B2(new_n524), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT119), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1051), .B(new_n392), .C1(new_n774), .C2(new_n1030), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1023), .B(new_n1278), .C1(new_n807), .C2(G107), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n458), .B2(new_n1036), .C1(new_n615), .C2(new_n1062), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1271), .A2(new_n1275), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1268), .B1(new_n1281), .B2(new_n815), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1267), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1257), .B2(new_n1166), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1264), .A2(new_n1285), .ZN(G381));
  OR2_X1    g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G384), .A2(new_n1287), .A3(G390), .A4(G381), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G387), .A2(new_n1288), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1089(.A1(new_n689), .A2(G213), .ZN(new_n1290));
  OR3_X1    g1090(.A1(G375), .A2(G378), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(G407), .A2(G213), .A3(new_n1291), .ZN(G409));
  INV_X1    g1092(.A(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1019), .A2(new_n1048), .A3(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G390), .B1(new_n1019), .B2(new_n1048), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT123), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1294), .A2(new_n1299), .A3(new_n1297), .A4(new_n1295), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1258), .A2(new_n1225), .A3(new_n1262), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT121), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1258), .A2(new_n1225), .A3(KEYINPUT121), .A4(new_n1262), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1256), .A2(new_n756), .A3(new_n1259), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1306), .A2(new_n1251), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G378), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G378), .B(new_n1252), .C1(new_n1254), .C2(new_n1260), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1134), .A2(new_n1142), .A3(new_n1124), .A4(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n709), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT60), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1263), .B1(new_n1143), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1319), .B2(new_n1285), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1321), .B(new_n1284), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1313), .A2(new_n1290), .A3(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(KEYINPUT63), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n689), .A2(G213), .A3(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT60), .B1(new_n1257), .B2(new_n1124), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1315), .B1(new_n1263), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1321), .B1(new_n1330), .B2(new_n1284), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1319), .A2(G384), .A3(new_n1285), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1326), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1334), .B1(new_n1313), .B2(new_n1290), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT122), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI22_X1  g1137(.A1(new_n1311), .A2(new_n1312), .B1(G213), .B2(new_n689), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT122), .B1(new_n1338), .B2(new_n1334), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1303), .A2(new_n1325), .A3(new_n1337), .A4(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1335), .B2(KEYINPUT61), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  OAI211_X1 g1143(.A(KEYINPUT124), .B(new_n1343), .C1(new_n1338), .C2(new_n1334), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT125), .ZN(new_n1346));
  AOI211_X1 g1146(.A(new_n1346), .B(KEYINPUT62), .C1(new_n1338), .C2(new_n1323), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT62), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT125), .B1(new_n1324), .B2(new_n1348), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1290), .A4(new_n1323), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(KEYINPUT126), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1345), .B1(new_n1350), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1340), .B1(new_n1353), .B2(new_n1354), .ZN(G405));
  NAND2_X1  g1155(.A1(new_n1354), .A2(KEYINPUT127), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT127), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1301), .A2(new_n1357), .A3(new_n1302), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1310), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1312), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1323), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1360), .A2(new_n1323), .ZN(new_n1363));
  OAI211_X1 g1163(.A(new_n1356), .B(new_n1358), .C1(new_n1362), .C2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1354), .A2(new_n1365), .A3(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(G402));
endmodule


