

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XNOR2_X1 U325 ( .A(KEYINPUT125), .B(n457), .ZN(n573) );
  XOR2_X1 U326 ( .A(n334), .B(n333), .Z(n532) );
  XOR2_X1 U327 ( .A(n374), .B(n399), .Z(n293) );
  XOR2_X1 U328 ( .A(n325), .B(KEYINPUT88), .Z(n294) );
  XOR2_X1 U329 ( .A(KEYINPUT93), .B(n467), .Z(n295) );
  XNOR2_X1 U330 ( .A(KEYINPUT25), .B(KEYINPUT94), .ZN(n468) );
  XNOR2_X1 U331 ( .A(n469), .B(n468), .ZN(n475) );
  XNOR2_X1 U332 ( .A(G176GAT), .B(G92GAT), .ZN(n323) );
  NOR2_X1 U333 ( .A1(n529), .A2(n476), .ZN(n477) );
  XNOR2_X1 U334 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n417) );
  XNOR2_X1 U335 ( .A(n418), .B(n417), .ZN(n419) );
  NOR2_X1 U336 ( .A1(n590), .A2(n492), .ZN(n493) );
  XOR2_X1 U337 ( .A(KEYINPUT41), .B(n583), .Z(n561) );
  XNOR2_X1 U338 ( .A(n498), .B(KEYINPUT38), .ZN(n507) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U340 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U341 ( .A(KEYINPUT72), .ZN(n296) );
  NAND2_X1 U342 ( .A1(G134GAT), .A2(n296), .ZN(n299) );
  INV_X1 U343 ( .A(G134GAT), .ZN(n297) );
  NAND2_X1 U344 ( .A1(n297), .A2(KEYINPUT72), .ZN(n298) );
  NAND2_X1 U345 ( .A1(n299), .A2(n298), .ZN(n354) );
  XOR2_X1 U346 ( .A(n354), .B(G162GAT), .Z(n303) );
  XOR2_X1 U347 ( .A(G127GAT), .B(KEYINPUT76), .Z(n301) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n445) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(n445), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n316) );
  XOR2_X1 U352 ( .A(G85GAT), .B(G148GAT), .Z(n305) );
  XNOR2_X1 U353 ( .A(G141GAT), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n307) );
  XNOR2_X1 U356 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(n309), .B(n308), .Z(n314) );
  XOR2_X1 U359 ( .A(KEYINPUT4), .B(KEYINPUT87), .Z(n311) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(n312), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U365 ( .A(KEYINPUT3), .B(KEYINPUT83), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT82), .B(G155GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(KEYINPUT2), .B(n319), .ZN(n436) );
  XOR2_X1 U369 ( .A(n320), .B(n436), .Z(n512) );
  INV_X1 U370 ( .A(n512), .ZN(n529) );
  XOR2_X1 U371 ( .A(KEYINPUT90), .B(G218GAT), .Z(n322) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n329) );
  XNOR2_X1 U374 ( .A(n323), .B(G64GAT), .ZN(n374) );
  XOR2_X1 U375 ( .A(G169GAT), .B(G8GAT), .Z(n399) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n293), .B(n324), .ZN(n325) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n326), .B(G211GAT), .ZN(n420) );
  XNOR2_X1 U380 ( .A(n420), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n294), .B(n327), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U383 ( .A(KEYINPUT19), .B(G190GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U386 ( .A(KEYINPUT18), .B(n332), .ZN(n453) );
  INV_X1 U387 ( .A(n453), .ZN(n333) );
  XOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .Z(n373) );
  XOR2_X1 U389 ( .A(G155GAT), .B(G71GAT), .Z(n336) );
  XNOR2_X1 U390 ( .A(G183GAT), .B(G127GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U392 ( .A(n373), .B(n337), .Z(n339) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(n340), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U396 ( .A(G15GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n341), .B(KEYINPUT67), .ZN(n401) );
  XNOR2_X1 U398 ( .A(n401), .B(G8GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT15), .B(G211GAT), .Z(n345) );
  XNOR2_X1 U401 ( .A(G22GAT), .B(G78GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n347) );
  XNOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(n349), .B(n348), .Z(n350) );
  XOR2_X1 U407 ( .A(n351), .B(n350), .Z(n494) );
  XOR2_X1 U408 ( .A(KEYINPUT11), .B(KEYINPUT71), .Z(n353) );
  XNOR2_X1 U409 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n364) );
  XOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .Z(n381) );
  XNOR2_X1 U412 ( .A(n381), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(G190GAT), .B(G106GAT), .Z(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n358) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U419 ( .A(G218GAT), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U420 ( .A(n421), .B(KEYINPUT73), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n370) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(G29GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n366), .B(KEYINPUT7), .ZN(n368) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(G50GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n396) );
  INV_X1 U428 ( .A(n396), .ZN(n369) );
  XOR2_X1 U429 ( .A(n370), .B(n369), .Z(n463) );
  XNOR2_X1 U430 ( .A(KEYINPUT36), .B(n463), .ZN(n590) );
  NOR2_X1 U431 ( .A1(n494), .A2(n590), .ZN(n372) );
  INV_X1 U432 ( .A(KEYINPUT45), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n387) );
  XOR2_X1 U434 ( .A(n374), .B(n373), .Z(n378) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G148GAT), .Z(n376) );
  XNOR2_X1 U437 ( .A(G106GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n431) );
  XNOR2_X1 U439 ( .A(n442), .B(n431), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n380) );
  XNOR2_X1 U442 ( .A(KEYINPUT31), .B(KEYINPUT70), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U444 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U445 ( .A1(G230GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n462) );
  INV_X1 U448 ( .A(n462), .ZN(n583) );
  NOR2_X1 U449 ( .A1(n387), .A2(n583), .ZN(n389) );
  INV_X1 U450 ( .A(KEYINPUT114), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n404) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n391) );
  NAND2_X1 U453 ( .A1(G229GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n392), .B(KEYINPUT29), .Z(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT65), .B(KEYINPUT68), .Z(n394) );
  XNOR2_X1 U457 ( .A(G113GAT), .B(G197GAT), .ZN(n393) );
  XOR2_X1 U458 ( .A(n394), .B(n393), .Z(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n403) );
  XOR2_X1 U462 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XNOR2_X1 U463 ( .A(n427), .B(n401), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT69), .ZN(n570) );
  NOR2_X1 U466 ( .A1(n404), .A2(n570), .ZN(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT115), .B(n405), .ZN(n414) );
  INV_X1 U468 ( .A(n494), .ZN(n587) );
  INV_X1 U469 ( .A(n406), .ZN(n579) );
  NAND2_X1 U470 ( .A1(n579), .A2(n561), .ZN(n407) );
  XOR2_X1 U471 ( .A(KEYINPUT46), .B(n407), .Z(n408) );
  NOR2_X1 U472 ( .A1(n587), .A2(n408), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n409), .B(KEYINPUT112), .ZN(n410) );
  NAND2_X1 U474 ( .A1(n410), .A2(n463), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n411), .B(KEYINPUT113), .ZN(n412) );
  XNOR2_X1 U476 ( .A(KEYINPUT47), .B(n412), .ZN(n413) );
  NAND2_X1 U477 ( .A1(n414), .A2(n413), .ZN(n416) );
  XNOR2_X1 U478 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n541) );
  NAND2_X1 U480 ( .A1(n532), .A2(n541), .ZN(n418) );
  NOR2_X1 U481 ( .A1(n529), .A2(n419), .ZN(n578) );
  XOR2_X1 U482 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n425) );
  XNOR2_X1 U486 ( .A(KEYINPUT81), .B(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U488 ( .A(n426), .B(KEYINPUT85), .Z(n429) );
  XNOR2_X1 U489 ( .A(G50GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U491 ( .A(n430), .B(KEYINPUT86), .Z(n433) );
  XNOR2_X1 U492 ( .A(n431), .B(KEYINPUT22), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n470) );
  NAND2_X1 U496 ( .A1(n578), .A2(n470), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n438), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U498 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(G134GAT), .Z(n444) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U504 ( .A(G169GAT), .B(n445), .Z(n447) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U507 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT77), .Z(n451) );
  XNOR2_X1 U509 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U511 ( .A(n453), .B(n452), .Z(n454) );
  XOR2_X1 U512 ( .A(n455), .B(n454), .Z(n520) );
  INV_X1 U513 ( .A(n520), .ZN(n544) );
  NAND2_X1 U514 ( .A1(n456), .A2(n544), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n573), .A2(n561), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT126), .B(KEYINPUT56), .Z(n459) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n483) );
  NAND2_X1 U519 ( .A1(n570), .A2(n462), .ZN(n497) );
  INV_X1 U520 ( .A(n463), .ZN(n574) );
  NOR2_X1 U521 ( .A1(n574), .A2(n494), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT16), .ZN(n480) );
  INV_X1 U523 ( .A(n532), .ZN(n516) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n516), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n512), .A2(n473), .ZN(n540) );
  XOR2_X1 U526 ( .A(KEYINPUT28), .B(n470), .Z(n537) );
  INV_X1 U527 ( .A(n537), .ZN(n543) );
  NAND2_X1 U528 ( .A1(n540), .A2(n543), .ZN(n465) );
  XOR2_X1 U529 ( .A(KEYINPUT91), .B(n465), .Z(n466) );
  NOR2_X1 U530 ( .A1(n544), .A2(n466), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n544), .A2(n532), .ZN(n467) );
  NAND2_X1 U532 ( .A1(n470), .A2(n295), .ZN(n469) );
  NOR2_X1 U533 ( .A1(n544), .A2(n470), .ZN(n472) );
  XNOR2_X1 U534 ( .A(KEYINPUT92), .B(KEYINPUT26), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(n577) );
  INV_X1 U536 ( .A(n577), .ZN(n559) );
  NOR2_X1 U537 ( .A1(n473), .A2(n559), .ZN(n474) );
  NOR2_X1 U538 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U539 ( .A1(n478), .A2(n477), .ZN(n492) );
  INV_X1 U540 ( .A(n492), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n510) );
  NOR2_X1 U542 ( .A1(n497), .A2(n510), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT95), .B(n481), .Z(n489) );
  NAND2_X1 U544 ( .A1(n489), .A2(n529), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U546 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  NAND2_X1 U547 ( .A1(n532), .A2(n489), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U550 ( .A1(n489), .A2(n544), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NAND2_X1 U553 ( .A1(n537), .A2(n489), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(KEYINPUT98), .ZN(n491) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U557 ( .A1(n494), .A2(n493), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n528) );
  NOR2_X1 U560 ( .A1(n528), .A2(n497), .ZN(n498) );
  NAND2_X1 U561 ( .A1(n507), .A2(n529), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U563 ( .A(G29GAT), .B(n501), .Z(G1328GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n532), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n504) );
  NAND2_X1 U568 ( .A1(n544), .A2(n507), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1330GAT) );
  XOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U572 ( .A1(n507), .A2(n537), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  NAND2_X1 U574 ( .A1(n561), .A2(n406), .ZN(n527) );
  NOR2_X1 U575 ( .A1(n510), .A2(n527), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT104), .B(n511), .Z(n522) );
  NOR2_X1 U577 ( .A1(n512), .A2(n522), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  XNOR2_X1 U581 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n516), .A2(n522), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(n519), .ZN(G1333GAT) );
  NOR2_X1 U585 ( .A1(n522), .A2(n520), .ZN(n521) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n543), .ZN(n526) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n524) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  XOR2_X1 U596 ( .A(G92GAT), .B(KEYINPUT111), .Z(n534) );
  NAND2_X1 U597 ( .A1(n536), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n544), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(n542), .Z(n558) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U607 ( .A1(n558), .A2(n545), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n570), .A2(n554), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n546), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U611 ( .A1(n554), .A2(n561), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT118), .Z(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT50), .Z(n552) );
  NAND2_X1 U616 ( .A1(n554), .A2(n587), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n553), .Z(G1342GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U620 ( .A1(n554), .A2(n574), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(G134GAT), .B(n557), .Z(G1343GAT) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n579), .A2(n567), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n587), .A2(n567), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT123), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n574), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n573), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n587), .A2(n573), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n589) );
  INV_X1 U645 ( .A(n589), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

