//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n196), .A2(KEYINPUT64), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n193), .A3(new_n195), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n192), .A3(G143), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n194), .B(G146), .C1(new_n203), .C2(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT82), .B(G224), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n219), .A2(KEYINPUT77), .A3(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT77), .B1(new_n219), .B2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n225), .B2(G104), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(KEYINPUT77), .A3(G107), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n223), .A4(new_n226), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G116), .B(G119), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT2), .B(G113), .Z(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n236), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G101), .C1(new_n222), .C2(new_n227), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n235), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  OR3_X1    g061(.A1(new_n247), .A2(KEYINPUT5), .A3(G119), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(G113), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n225), .B2(G104), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n225), .A2(G104), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n219), .A2(KEYINPUT78), .A3(G107), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n241), .A3(new_n234), .A4(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G122), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n245), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(KEYINPUT8), .ZN(new_n259));
  INV_X1    g073(.A(new_n256), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n249), .A2(new_n241), .B1(new_n234), .B2(new_n255), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n202), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n211), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n218), .A2(new_n258), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n256), .ZN(new_n267));
  INV_X1    g081(.A(new_n257), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n258), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n245), .A2(new_n256), .A3(new_n257), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n257), .B1(new_n245), .B2(new_n256), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n267), .A2(new_n273), .A3(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n270), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n212), .B(new_n216), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n266), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n187), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n282), .A2(KEYINPUT83), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n258), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT81), .B1(new_n272), .B2(new_n273), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n288), .B2(new_n270), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n284), .A2(new_n187), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n289), .A2(new_n266), .A3(new_n290), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n283), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n235), .A2(new_n297), .A3(new_n244), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT11), .ZN(new_n299));
  INV_X1    g113(.A(G134), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(G137), .ZN(new_n301));
  INV_X1    g115(.A(G137), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT11), .A3(G134), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(G137), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G131), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n301), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n234), .A2(new_n208), .A3(new_n255), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n234), .A2(new_n255), .A3(new_n208), .A4(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n298), .A2(new_n309), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n308), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n315), .A2(KEYINPUT79), .ZN(new_n316));
  INV_X1    g130(.A(new_n310), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n208), .B1(new_n234), .B2(new_n255), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT12), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n215), .A2(G227), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n316), .B(new_n324), .C1(new_n317), .C2(new_n318), .ZN(new_n325));
  AND4_X1   g139(.A1(new_n314), .A2(new_n320), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n235), .A2(new_n297), .A3(new_n244), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n312), .A2(new_n313), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n327), .B(new_n315), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n298), .A2(new_n312), .A3(new_n313), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(new_n315), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n314), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n323), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(G469), .A3(G902), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n315), .B1(new_n328), .B2(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT80), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n330), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n314), .A2(new_n323), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n320), .A2(new_n314), .A3(new_n325), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n335), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n344), .A3(G469), .ZN(new_n345));
  INV_X1    g159(.A(G469), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(new_n265), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n293), .B(new_n296), .C1(new_n337), .C2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n219), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n210), .A2(G140), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT16), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(new_n354), .A3(KEYINPUT69), .A4(G125), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n192), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n356), .A2(new_n358), .A3(G146), .A4(new_n360), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(KEYINPUT70), .A3(new_n192), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  AND2_X1   g182(.A1(KEYINPUT85), .A2(G143), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT85), .A2(G143), .ZN(new_n370));
  OAI211_X1 g184(.A(G214), .B(new_n368), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n215), .A3(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(KEYINPUT85), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n307), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT17), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n368), .A2(G214), .B1(KEYINPUT85), .B2(G143), .ZN(new_n378));
  INV_X1    g192(.A(new_n373), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT85), .B(G143), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n307), .ZN(new_n382));
  INV_X1    g196(.A(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n367), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n355), .A2(new_n357), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n192), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n355), .A2(new_n357), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n376), .A2(KEYINPUT18), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n371), .B(new_n375), .C1(new_n392), .C2(new_n307), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT87), .B(new_n391), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n381), .B(new_n398), .C1(new_n392), .C2(new_n307), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT87), .B1(new_n401), .B2(new_n391), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n352), .B(new_n386), .C1(new_n397), .C2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n382), .A2(new_n383), .ZN(new_n407));
  INV_X1    g221(.A(new_n364), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n387), .A2(KEYINPUT88), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n411), .B2(new_n192), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n406), .A2(new_n396), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n403), .B1(new_n413), .B2(new_n352), .ZN(new_n414));
  INV_X1    g228(.A(G475), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n265), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n414), .A2(new_n418), .A3(new_n415), .A4(new_n265), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n215), .A2(G952), .ZN(new_n421));
  NAND2_X1  g235(.A1(G234), .A2(G237), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT90), .Z(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(G902), .A3(G953), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G116), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(G107), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT89), .ZN(new_n435));
  XNOR2_X1  g249(.A(G128), .B(G143), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n300), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n194), .A2(G128), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n438), .B(G134), .C1(KEYINPUT13), .C2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n436), .B(new_n300), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n247), .A2(KEYINPUT14), .A3(G122), .ZN(new_n443));
  INV_X1    g257(.A(new_n433), .ZN(new_n444));
  OAI211_X1 g258(.A(G107), .B(new_n443), .C1(new_n444), .C2(KEYINPUT14), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n442), .B(new_n445), .C1(G107), .C2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G217), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n295), .A2(new_n448), .A3(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(new_n446), .A3(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n432), .B1(new_n453), .B2(new_n265), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n441), .A2(new_n446), .A3(new_n449), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n441), .B2(new_n446), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n265), .B(new_n432), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n386), .B1(new_n397), .B2(new_n402), .ZN(new_n460));
  INV_X1    g274(.A(new_n352), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n403), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n265), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G475), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n420), .A2(new_n429), .A3(new_n459), .A4(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n292), .A2(new_n350), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n468));
  INV_X1    g282(.A(G472), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n242), .B(KEYINPUT66), .ZN(new_n470));
  INV_X1    g284(.A(new_n304), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n300), .A2(G137), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n208), .A2(new_n308), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n309), .B2(new_n201), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n242), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n315), .A2(new_n200), .A3(new_n191), .A4(new_n199), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n474), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n368), .A2(G210), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n233), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n470), .A2(new_n475), .ZN(new_n488));
  AND4_X1   g302(.A1(KEYINPUT29), .A2(new_n482), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n475), .A2(new_n242), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n486), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n242), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n495), .A2(KEYINPUT65), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(KEYINPUT65), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n475), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n480), .A2(KEYINPUT65), .A3(new_n495), .A4(new_n474), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n470), .A2(new_n475), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n500), .A2(new_n501), .A3(new_n487), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n491), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n469), .B1(new_n490), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n506), .B2(new_n242), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n507), .B2(new_n487), .ZN(new_n508));
  NOR4_X1   g322(.A1(new_n500), .A2(KEYINPUT31), .A3(new_n501), .A4(new_n486), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n487), .B1(new_n482), .B2(new_n492), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G472), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT32), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n487), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n516));
  INV_X1    g330(.A(new_n510), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n507), .A2(new_n505), .A3(new_n487), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n512), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n504), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G110), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G119), .B(G128), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT23), .B1(new_n203), .B2(G119), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n203), .A2(G119), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT68), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n532));
  OAI211_X1 g346(.A(G119), .B(new_n203), .C1(new_n532), .C2(KEYINPUT23), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G110), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n365), .A2(new_n528), .A3(new_n535), .A4(new_n366), .ZN(new_n536));
  NOR2_X1   g350(.A1(KEYINPUT71), .A2(G110), .ZN(new_n537));
  AND2_X1   g351(.A1(KEYINPUT71), .A2(G110), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n364), .B(new_n388), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT72), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n536), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n545), .B1(new_n536), .B2(new_n541), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n265), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n448), .B1(G234), .B2(new_n265), .ZN(new_n549));
  OR3_X1    g363(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT75), .B1(new_n548), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n536), .A2(new_n541), .ZN(new_n553));
  INV_X1    g367(.A(new_n545), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n536), .A2(new_n541), .A3(new_n545), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT73), .B1(new_n557), .B2(KEYINPUT25), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT25), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT25), .B(new_n265), .C1(new_n546), .C2(new_n547), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT73), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n548), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n558), .A2(new_n560), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n552), .B1(new_n549), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n468), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n504), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n511), .A2(KEYINPUT32), .A3(new_n513), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n520), .B1(new_n519), .B2(new_n512), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT76), .A3(new_n567), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n467), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  XNOR2_X1  g390(.A(new_n409), .B(KEYINPUT19), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n364), .B(new_n407), .C1(new_n577), .C2(G146), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n397), .B2(new_n402), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n461), .ZN(new_n580));
  AOI21_X1  g394(.A(G475), .B1(new_n580), .B2(new_n403), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n418), .B1(new_n581), .B2(new_n265), .ZN(new_n582));
  AND4_X1   g396(.A1(new_n418), .A2(new_n414), .A3(new_n415), .A4(new_n265), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n465), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT33), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n455), .B2(new_n456), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n451), .A2(KEYINPUT33), .A3(new_n452), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n430), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n430), .B(new_n265), .C1(new_n455), .C2(new_n456), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n430), .A2(new_n265), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n278), .A2(new_n280), .ZN(new_n594));
  INV_X1    g408(.A(new_n266), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n282), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n282), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n597), .B(new_n266), .C1(new_n278), .C2(new_n280), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n293), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n593), .A2(new_n599), .A3(new_n428), .ZN(new_n600));
  INV_X1    g414(.A(new_n296), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n323), .B1(new_n340), .B2(new_n314), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n346), .B(new_n265), .C1(new_n602), .C2(new_n326), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n340), .A2(new_n341), .B1(new_n335), .B2(new_n343), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n347), .B1(new_n604), .B2(G469), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT91), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n519), .B(new_n265), .C1(new_n607), .C2(new_n469), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT91), .B(G472), .C1(new_n511), .C2(G902), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n567), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(new_n293), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n594), .A2(new_n282), .A3(new_n595), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n597), .B1(new_n289), .B2(new_n266), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n419), .A2(KEYINPUT92), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n581), .A2(new_n619), .A3(new_n418), .A4(new_n265), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n620), .A3(new_n417), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n465), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n459), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n610), .A2(new_n429), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n350), .A2(new_n466), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n281), .A2(new_n284), .ZN(new_n629));
  INV_X1    g443(.A(new_n291), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n608), .A2(new_n609), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n566), .A2(new_n549), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n553), .B1(KEYINPUT36), .B2(new_n545), .ZN(new_n634));
  INV_X1    g448(.A(new_n549), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n545), .A2(KEYINPUT36), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n536), .A3(new_n541), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n634), .A2(new_n265), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT93), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n627), .A2(new_n631), .A3(new_n632), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(new_n459), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n424), .B(KEYINPUT94), .Z(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n425), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n646), .A2(new_n621), .A3(new_n465), .A4(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n640), .B1(new_n566), .B2(new_n549), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n599), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n654), .A3(new_n573), .A4(new_n606), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  OAI21_X1  g470(.A(new_n487), .B1(new_n500), .B2(new_n501), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n501), .A2(new_n487), .ZN(new_n659));
  AOI211_X1 g473(.A(G902), .B(new_n658), .C1(new_n488), .C2(new_n659), .ZN(new_n660));
  OAI22_X1  g474(.A1(new_n571), .A2(new_n572), .B1(new_n469), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT96), .Z(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n292), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n584), .A2(new_n646), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n650), .B(KEYINPUT39), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n606), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n653), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n293), .B1(new_n670), .B2(new_n671), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n663), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n194), .ZN(G45));
  AOI21_X1  g490(.A(new_n415), .B1(new_n463), .B2(new_n265), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n417), .B2(new_n419), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n586), .A2(new_n587), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G478), .ZN(new_n680));
  INV_X1    g494(.A(new_n591), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n589), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n678), .A2(new_n682), .A3(new_n650), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n654), .A2(new_n683), .A3(new_n573), .A4(new_n606), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT97), .B(G146), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  NOR2_X1   g500(.A1(new_n522), .A2(new_n568), .ZN(new_n687));
  OAI21_X1  g501(.A(G469), .B1(new_n336), .B2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n296), .A3(new_n603), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n600), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n599), .A2(new_n689), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n687), .A2(new_n429), .A3(new_n623), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n522), .A2(new_n466), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n642), .A3(new_n694), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  OAI21_X1  g513(.A(G472), .B1(new_n511), .B2(G902), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n512), .B(KEYINPUT98), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n516), .A2(new_n518), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n487), .B1(new_n482), .B2(new_n488), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n568), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n666), .A2(new_n599), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n429), .A4(new_n690), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT99), .B(G122), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G24));
  NOR2_X1   g524(.A1(new_n705), .A2(new_n653), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n694), .A3(new_n683), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n293), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n603), .A2(new_n605), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n296), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n292), .A2(KEYINPUT100), .A3(new_n293), .A4(new_n606), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n687), .A3(new_n683), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n584), .A2(new_n592), .A3(new_n651), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n522), .B2(new_n568), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n722), .B1(new_n718), .B2(new_n719), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n307), .ZN(G33));
  AND3_X1   g546(.A1(new_n720), .A2(new_n687), .A3(new_n652), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n300), .ZN(G36));
  OAI21_X1  g548(.A(G469), .B1(new_n604), .B2(KEYINPUT45), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT102), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n604), .A2(KEYINPUT45), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n347), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n742), .A3(KEYINPUT46), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n741), .A3(new_n603), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n296), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n667), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n678), .A2(new_n592), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n632), .A3(new_n653), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n715), .B1(new_n752), .B2(KEYINPUT44), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n746), .B(new_n753), .C1(KEYINPUT44), .C2(new_n752), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  NOR3_X1   g569(.A1(new_n573), .A2(new_n715), .A3(new_n567), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n296), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT47), .B1(new_n744), .B2(new_n296), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n683), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n688), .A2(new_n603), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n747), .B(new_n665), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n761), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n567), .A2(new_n293), .A3(new_n296), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT105), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(new_n663), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n751), .A2(new_n647), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n689), .A2(new_n293), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n665), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(new_n770), .A3(new_n706), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n774), .A2(new_n776), .A3(KEYINPUT115), .A4(new_n775), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n779), .B(new_n780), .C1(new_n775), .C2(new_n773), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n715), .A2(new_n689), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n768), .A2(new_n711), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT116), .Z(new_n784));
  NOR2_X1   g598(.A1(new_n757), .A2(new_n758), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n762), .A2(new_n601), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n715), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n768), .A2(new_n706), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n568), .A2(new_n424), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n663), .A2(new_n782), .A3(new_n790), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(new_n584), .A3(new_n592), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n781), .A2(new_n789), .A3(KEYINPUT51), .A4(new_n792), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n791), .A2(new_n593), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n421), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n678), .A2(new_n646), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n428), .B1(new_n593), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n610), .A2(new_n800), .A3(new_n631), .A4(new_n293), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n575), .A2(new_n801), .A3(new_n643), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT106), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n575), .A2(new_n801), .A3(KEYINPUT106), .A4(new_n643), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n733), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n691), .A2(new_n695), .A3(new_n708), .A4(new_n698), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n723), .B2(new_n730), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n593), .B(new_n705), .C1(new_n718), .C2(new_n719), .ZN(new_n809));
  INV_X1    g623(.A(new_n715), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n573), .A3(new_n606), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n646), .A3(new_n622), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n642), .B(new_n651), .C1(new_n809), .C2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n806), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n642), .A2(new_n617), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n522), .A3(new_n717), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n548), .A2(new_n563), .A3(new_n564), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n563), .B1(new_n548), .B2(new_n564), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n561), .B(new_n559), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n635), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n700), .B(new_n704), .C1(new_n822), .C2(new_n640), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n724), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n817), .A2(new_n652), .B1(new_n824), .B2(new_n694), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n651), .A2(KEYINPUT107), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n651), .A2(KEYINPUT107), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n296), .A2(new_n716), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n707), .A2(new_n828), .A3(new_n653), .A4(new_n661), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n825), .A2(KEYINPUT109), .A3(new_n684), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n655), .A3(new_n684), .A4(new_n712), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n830), .A2(KEYINPUT52), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n830), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n815), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n833), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT52), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(KEYINPUT110), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n814), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n831), .A2(new_n838), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT108), .B1(new_n835), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(KEYINPUT108), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n806), .A2(new_n813), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n808), .A2(KEYINPUT111), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n843), .B1(new_n808), .B2(KEYINPUT111), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n844), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n788), .A2(new_n694), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n849), .A2(new_n843), .A3(new_n814), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n844), .A2(new_n853), .A3(new_n860), .A4(new_n845), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n856), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n725), .A2(new_n727), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n768), .A2(new_n863), .A3(new_n782), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n798), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n767), .B1(new_n867), .B2(new_n868), .ZN(G75));
  AOI21_X1  g683(.A(new_n265), .B1(new_n844), .B2(new_n853), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(G210), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n278), .B(KEYINPUT118), .Z(new_n872));
  XNOR2_X1  g686(.A(new_n279), .B(KEYINPUT55), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(KEYINPUT56), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n871), .A2(new_n876), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n215), .A2(G952), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G51));
  NAND2_X1  g694(.A1(new_n348), .A2(KEYINPUT57), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n348), .A2(KEYINPUT57), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n844), .A2(new_n845), .A3(new_n853), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n845), .B1(new_n844), .B2(new_n853), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n602), .B2(new_n326), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n870), .A2(new_n737), .A3(new_n736), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(G54));
  NAND3_X1  g702(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(new_n414), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n879), .ZN(G60));
  NAND3_X1  g705(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n892));
  XNOR2_X1  g706(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n681), .B(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n679), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  INV_X1    g712(.A(new_n679), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n895), .C1(new_n883), .C2(new_n884), .ZN(new_n900));
  INV_X1    g714(.A(new_n879), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n892), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(new_n844), .A2(new_n853), .ZN(new_n908));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT60), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n634), .A2(new_n637), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n901), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT61), .B1(new_n914), .B2(KEYINPUT122), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n556), .A3(new_n555), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n916), .B(new_n901), .C1(new_n913), .C2(new_n911), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n915), .B(new_n917), .ZN(G66));
  AND2_X1   g732(.A1(new_n804), .A2(new_n805), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(new_n807), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n215), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT123), .Z(new_n922));
  INV_X1    g736(.A(new_n214), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n923), .B2(new_n426), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n872), .B1(G898), .B2(new_n215), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  AOI21_X1  g741(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n506), .B(new_n577), .ZN(new_n929));
  XOR2_X1   g743(.A(KEYINPUT125), .B(G900), .Z(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n929), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n825), .A2(new_n684), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n675), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n675), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n569), .A2(new_n574), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n593), .B2(new_n799), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n670), .A3(new_n810), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n937), .A2(new_n754), .A3(new_n759), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n932), .B1(new_n941), .B2(new_n215), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n928), .ZN(new_n943));
  INV_X1    g757(.A(new_n733), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n754), .A2(new_n944), .A3(new_n759), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n746), .A2(new_n707), .A3(new_n863), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n731), .A2(new_n934), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n215), .B(new_n932), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT124), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n949), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  NOR4_X1   g766(.A1(new_n951), .A2(new_n942), .A3(new_n952), .A4(new_n928), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n931), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(new_n931), .C1(new_n950), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OR2_X1    g774(.A1(new_n945), .A2(new_n948), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n920), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n879), .B1(new_n962), .B2(new_n502), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n941), .B2(new_n920), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n658), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n657), .A2(new_n960), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n502), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n857), .A2(new_n858), .A3(new_n969), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n963), .A2(new_n966), .A3(new_n967), .A4(new_n970), .ZN(G57));
endmodule


