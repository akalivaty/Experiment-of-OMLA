//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT69), .A2(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT69), .A2(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G119), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT5), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G113), .ZN(new_n198));
  INV_X1    g012(.A(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT5), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n208), .A3(new_n204), .A4(G104), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n204), .A2(G104), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n207), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n194), .A3(new_n196), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n217), .B2(new_n210), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n202), .A2(new_n212), .A3(new_n215), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n202), .A2(new_n215), .B1(new_n212), .B2(new_n218), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n191), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G224), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT86), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G125), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT0), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT64), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n234), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g055(.A(G143), .B(G146), .ZN(new_n242));
  INV_X1    g056(.A(new_n234), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n237), .A2(new_n239), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n241), .A3(new_n233), .A4(new_n234), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n228), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n233), .A2(new_n250), .A3(G128), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n230), .B(new_n232), .C1(KEYINPUT1), .C2(new_n236), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G125), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n227), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n227), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n248), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n222), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT69), .A2(G116), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT69), .A2(G116), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n262), .A2(new_n263), .A3(new_n195), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n213), .B1(new_n264), .B2(new_n199), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n215), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n206), .A2(new_n211), .ZN(new_n268));
  INV_X1    g082(.A(new_n209), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n267), .B(G101), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n210), .B1(new_n205), .B2(KEYINPUT3), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n207), .B1(new_n272), .B2(new_n209), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n266), .B(new_n270), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT85), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n273), .A2(new_n267), .B1(new_n265), .B2(new_n215), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(KEYINPUT85), .A3(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n276), .A2(new_n280), .A3(new_n189), .A4(new_n219), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n222), .B(KEYINPUT89), .C1(new_n256), .C2(new_n258), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n261), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n189), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n219), .B1(new_n274), .B2(new_n275), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT85), .B1(new_n278), .B2(new_n279), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT6), .A3(new_n281), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n248), .A2(new_n254), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(new_n225), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT87), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT87), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n290), .A2(new_n297), .A3(new_n294), .A4(new_n292), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n285), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT90), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n188), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI211_X1 g115(.A(KEYINPUT90), .B(new_n285), .C1(new_n296), .C2(new_n298), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n188), .B(new_n285), .C1(new_n296), .C2(new_n298), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G475), .ZN(new_n306));
  XNOR2_X1  g120(.A(G125), .B(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n308));
  OR3_X1    g122(.A1(new_n228), .A2(KEYINPUT16), .A3(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(G146), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(G146), .B1(new_n308), .B2(new_n309), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT67), .B(G131), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(KEYINPUT71), .A2(G237), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT71), .A2(G237), .ZN(new_n317));
  AOI21_X1  g131(.A(G953), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G143), .B1(new_n318), .B2(G214), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT71), .A2(G237), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT71), .A2(G237), .ZN(new_n321));
  OAI211_X1 g135(.A(G214), .B(new_n223), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(new_n231), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n315), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT91), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n231), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT71), .B(G237), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(G143), .A3(G214), .A4(new_n223), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n315), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n313), .B1(new_n332), .B2(KEYINPUT17), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n328), .A3(new_n314), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n325), .A2(new_n334), .A3(new_n331), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT92), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n330), .B1(new_n329), .B2(new_n315), .ZN(new_n338));
  AOI211_X1 g152(.A(KEYINPUT91), .B(new_n314), .C1(new_n326), .C2(new_n328), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n334), .A4(new_n335), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n216), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n329), .A2(KEYINPUT18), .A3(G131), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n329), .B1(KEYINPUT18), .B2(G131), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n307), .B(G146), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n343), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(new_n345), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g169(.A(KEYINPUT93), .B(new_n345), .C1(new_n343), .C2(new_n350), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n306), .B1(new_n357), .B2(new_n284), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n307), .B(KEYINPUT19), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n360), .A2(new_n229), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n311), .B(new_n361), .C1(new_n340), .C2(new_n335), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n354), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n359), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  AOI211_X1 g181(.A(KEYINPUT20), .B(new_n367), .C1(new_n351), .C2(new_n363), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n358), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(G234), .A2(G237), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G952), .A3(new_n223), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT21), .B(G898), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n372), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G478), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(KEYINPUT15), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n381), .A2(new_n382), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G134), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n236), .A2(G143), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n231), .A2(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n236), .A2(G143), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT13), .ZN(new_n391));
  XNOR2_X1  g205(.A(G128), .B(G143), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT66), .B(G134), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n388), .A2(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n192), .A2(G122), .A3(new_n193), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n395), .A2(new_n204), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n204), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n394), .B(KEYINPUT94), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n398), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n392), .B(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n192), .A2(new_n408), .A3(G122), .A4(new_n193), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n410), .B1(G116), .B2(new_n396), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n395), .A2(new_n413), .A3(KEYINPUT14), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n395), .B2(KEYINPUT14), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n407), .B1(new_n416), .B2(G107), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n384), .B1(new_n404), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(G107), .ZN(new_n419));
  INV_X1    g233(.A(new_n407), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n402), .B2(new_n403), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n383), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n380), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AOI211_X1 g241(.A(KEYINPUT97), .B(G902), .C1(new_n418), .C2(new_n422), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n380), .B1(new_n430), .B2(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n370), .A2(new_n378), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n305), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G472), .A2(G902), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT73), .Z(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n385), .A2(KEYINPUT66), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G134), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n444), .A3(G137), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n385), .A2(G137), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n441), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n444), .ZN(new_n449));
  INV_X1    g263(.A(G137), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT11), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n441), .B1(new_n393), .B2(G137), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n393), .B2(G137), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n314), .B(new_n453), .C1(new_n454), .C2(new_n441), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n245), .A2(KEYINPUT70), .A3(new_n247), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT70), .B1(new_n245), .B2(new_n247), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n450), .A2(G134), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n393), .A2(G137), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n253), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n440), .B1(new_n459), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n245), .A2(new_n247), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n468), .A2(new_n440), .A3(new_n465), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n266), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n266), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n459), .A2(new_n471), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n318), .A2(G210), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT27), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G101), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n470), .A2(new_n477), .A3(KEYINPUT72), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT72), .B1(new_n470), .B2(new_n477), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT31), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n472), .A2(new_n476), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT70), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n484), .A2(new_n485), .B1(new_n455), .B2(new_n452), .ZN(new_n486));
  INV_X1    g300(.A(new_n465), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT30), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n468), .A2(new_n440), .A3(new_n465), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n482), .B1(new_n490), .B2(new_n266), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n480), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n468), .A2(new_n465), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n266), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n459), .A2(KEYINPUT28), .A3(new_n471), .A4(new_n465), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n475), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n474), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n439), .B1(new_n481), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n471), .B1(new_n488), .B2(new_n489), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n482), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n470), .A2(new_n477), .A3(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT31), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n491), .A2(new_n480), .B1(new_n500), .B2(new_n498), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n438), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n500), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n266), .B1(new_n486), .B2(new_n487), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n494), .A2(new_n517), .A3(new_n497), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n284), .B1(new_n519), .B2(KEYINPUT75), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(KEYINPUT76), .A3(new_n284), .A4(new_n520), .ZN(new_n525));
  INV_X1    g339(.A(new_n472), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n500), .B1(new_n507), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n516), .C1(new_n500), .C2(new_n498), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n504), .A2(new_n514), .B1(G472), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n382), .B1(G234), .B2(new_n284), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT22), .B(G137), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n307), .A2(new_n229), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n310), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT23), .A2(G119), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(G128), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n236), .A2(KEYINPUT77), .A3(KEYINPUT23), .A4(G119), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G110), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n195), .A2(G128), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n236), .A2(G119), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT78), .B1(new_n544), .B2(KEYINPUT23), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n542), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n546), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT80), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n537), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n550), .A2(new_n551), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n311), .B2(new_n312), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT79), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(G110), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n559), .A3(G110), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n535), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n555), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n536), .B(new_n310), .C1(new_n566), .C2(new_n553), .ZN(new_n567));
  INV_X1    g381(.A(new_n563), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n313), .B(new_n557), .C1(new_n568), .C2(new_n561), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n569), .A3(new_n534), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT81), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT81), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  AOI211_X1 g388(.A(G902), .B(new_n531), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n531), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n570), .A3(new_n284), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT25), .A4(new_n284), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT82), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT82), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n572), .A2(new_n574), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n531), .A2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G469), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n223), .A2(G227), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n212), .A2(new_n218), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n253), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT84), .B1(new_n596), .B2(KEYINPUT10), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT84), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n598), .B(new_n599), .C1(new_n595), .C2(new_n253), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(KEYINPUT10), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n278), .B(new_n270), .C1(new_n457), .C2(new_n458), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n456), .ZN(new_n605));
  INV_X1    g419(.A(new_n456), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n601), .A2(new_n606), .A3(new_n602), .A4(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n594), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n212), .A2(new_n218), .B1(new_n251), .B2(new_n252), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n456), .B1(new_n596), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n456), .B(KEYINPUT12), .C1(new_n596), .C2(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n607), .A2(new_n594), .A3(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n590), .B(new_n284), .C1(new_n608), .C2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n607), .A2(new_n594), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n605), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n607), .A2(new_n614), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n593), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(G469), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(G469), .A2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n530), .A2(new_n589), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n436), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  NOR2_X1   g442(.A1(new_n379), .A2(G902), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n404), .A2(new_n417), .A3(new_n384), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n419), .A2(new_n420), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n402), .A2(new_n403), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n383), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT33), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n418), .B(new_n422), .C1(KEYINPUT101), .C2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n629), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  INV_X1    g456(.A(new_n427), .ZN(new_n643));
  INV_X1    g457(.A(new_n428), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n379), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n418), .A2(KEYINPUT101), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n646), .B(KEYINPUT33), .C1(new_n630), .C2(new_n633), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n629), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n642), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n378), .C1(new_n358), .C2(new_n369), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n299), .B2(new_n187), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n435), .B1(new_n299), .B2(new_n187), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n435), .A2(KEYINPUT100), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n304), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n660), .A3(KEYINPUT103), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n655), .A2(new_n656), .B1(new_n304), .B2(new_n658), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n652), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(G902), .B1(new_n510), .B2(new_n511), .ZN(new_n666));
  INV_X1    g480(.A(G472), .ZN(new_n667));
  OR3_X1    g481(.A1(new_n666), .A2(KEYINPUT99), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT99), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n503), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n589), .ZN(new_n671));
  INV_X1    g485(.A(new_n624), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n617), .A2(new_n605), .B1(new_n619), .B2(new_n593), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n672), .B1(new_n674), .B2(new_n616), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n665), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(new_n432), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n378), .A2(new_n660), .A3(new_n370), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT35), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  OAI22_X1  g499(.A1(new_n556), .A2(new_n564), .B1(KEYINPUT36), .B2(new_n535), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n569), .A2(new_n567), .A3(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n686), .A2(new_n688), .A3(new_n586), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n581), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n675), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n670), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n436), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT37), .B(G110), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT104), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G12));
  NOR3_X1   g511(.A1(new_n530), .A2(new_n625), .A3(new_n690), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G953), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n373), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n701), .B1(new_n373), .B2(new_n700), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n372), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n358), .A2(new_n369), .A3(new_n432), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n660), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n529), .A2(G472), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT32), .B1(new_n503), .B2(KEYINPUT74), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n512), .A2(new_n513), .A3(new_n505), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n675), .A3(new_n660), .A4(new_n691), .ZN(new_n713));
  INV_X1    g527(.A(new_n706), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XNOR2_X1  g531(.A(new_n305), .B(KEYINPUT38), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n704), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n675), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n434), .B(new_n690), .C1(new_n722), .C2(KEYINPUT40), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(KEYINPUT40), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n370), .A2(new_n432), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n518), .A2(new_n472), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n500), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n508), .A2(new_n509), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n284), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n710), .B2(new_n711), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n719), .A2(new_n724), .A3(new_n725), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  OAI211_X1 g549(.A(new_n651), .B(new_n704), .C1(new_n358), .C2(new_n369), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n713), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n229), .ZN(G48));
  OR2_X1    g552(.A1(new_n608), .A2(new_n615), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n284), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n624), .A3(new_n616), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n530), .A2(new_n589), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n665), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND2_X1  g560(.A1(new_n682), .A2(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR3_X1   g562(.A1(new_n530), .A2(new_n433), .A3(new_n690), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n742), .B1(new_n657), .B2(new_n659), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT109), .B(G119), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G21));
  INV_X1    g567(.A(new_n742), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n378), .A2(new_n725), .A3(new_n660), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n284), .B1(new_n481), .B2(new_n502), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(G472), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n666), .B2(new_n667), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n575), .A2(new_n581), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n494), .A2(new_n497), .A3(new_n518), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n491), .A2(new_n480), .B1(new_n500), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n438), .B1(new_n510), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n764), .B1(new_n758), .B2(new_n759), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT111), .B1(new_n769), .B2(new_n761), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n755), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  INV_X1    g586(.A(new_n736), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n750), .A2(new_n691), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n503), .A2(KEYINPUT32), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n512), .A2(new_n505), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n778), .B1(G472), .B2(new_n529), .ZN(new_n779));
  INV_X1    g593(.A(new_n761), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n779), .A2(new_n780), .A3(new_n736), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n675), .B(new_n656), .C1(new_n301), .C2(new_n302), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n776), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n736), .A2(KEYINPUT42), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n712), .A2(new_n785), .A3(new_n671), .A4(new_n783), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT112), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n777), .A2(new_n778), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n709), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n773), .A3(new_n761), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT42), .B1(new_n790), .B2(new_n782), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n530), .A2(new_n589), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n783), .A3(new_n785), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(G131), .Z(G33));
  NAND4_X1  g611(.A1(new_n712), .A2(new_n783), .A3(new_n671), .A4(new_n706), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  NAND2_X1  g613(.A1(new_n618), .A2(new_n620), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n590), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n622), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT46), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT113), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n616), .B1(new_n804), .B2(KEYINPUT46), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n624), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n656), .B1(new_n301), .B2(new_n302), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n721), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n370), .A2(new_n651), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT43), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n670), .A3(new_n691), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n813), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n814), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n450), .ZN(G39));
  NAND4_X1  g638(.A1(new_n530), .A2(new_n773), .A3(new_n812), .A4(new_n589), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n809), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(G140), .Z(G42));
  NOR2_X1   g644(.A1(new_n817), .A2(new_n372), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n768), .A2(new_n770), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n435), .A3(new_n718), .A4(new_n754), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT50), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n754), .A3(new_n812), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n690), .B(new_n764), .C1(new_n758), .C2(new_n759), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n812), .A2(new_n754), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n840), .A2(new_n733), .A3(new_n372), .A4(new_n589), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n370), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n651), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n835), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n833), .A2(new_n812), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n826), .A2(new_n828), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n741), .A2(new_n616), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n624), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n836), .A2(new_n780), .A3(new_n779), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT48), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(KEYINPUT120), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n833), .A2(new_n750), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n843), .A2(new_n651), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n223), .C1(new_n842), .C2(new_n858), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n854), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n849), .B(KEYINPUT119), .Z(new_n862));
  OAI21_X1  g676(.A(new_n846), .B1(new_n847), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n845), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n581), .A2(new_n689), .A3(new_n705), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n623), .A3(new_n624), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT116), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n675), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n733), .A2(new_n871), .A3(new_n660), .A4(new_n725), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n774), .B(new_n872), .C1(new_n713), .C2(new_n736), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n716), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n716), .A2(new_n874), .A3(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  MUX2_X1   g693(.A(new_n879), .B(new_n878), .S(KEYINPUT117), .Z(new_n880));
  NAND4_X1  g694(.A1(new_n783), .A2(new_n769), .A3(new_n773), .A4(new_n691), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n837), .A2(new_n883), .A3(new_n773), .A4(new_n783), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n366), .A2(new_n368), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n705), .B1(new_n429), .B2(new_n431), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n353), .A2(new_n354), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT93), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n353), .A2(new_n352), .A3(new_n354), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(G902), .B1(new_n891), .B2(new_n351), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n886), .B(new_n887), .C1(new_n892), .C2(new_n306), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n811), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n712), .A3(new_n675), .A4(new_n691), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(new_n798), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n858), .B1(new_n843), .B2(new_n432), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n305), .A2(new_n435), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n677), .A3(new_n898), .A4(new_n378), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n436), .B1(new_n626), .B2(new_n693), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n885), .A2(new_n896), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n771), .A2(new_n744), .A3(new_n747), .A4(new_n751), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n796), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  INV_X1    g720(.A(new_n796), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n716), .A2(new_n874), .A3(KEYINPUT52), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT52), .B1(new_n716), .B2(new_n874), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n880), .A2(new_n905), .B1(KEYINPUT53), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n791), .A2(new_n793), .A3(KEYINPUT53), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n901), .A2(new_n902), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n913), .B(new_n915), .C1(new_n879), .C2(KEYINPUT117), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n918), .B(KEYINPUT53), .C1(new_n879), .C2(new_n903), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT118), .B1(new_n910), .B2(new_n904), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n916), .B(new_n917), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n865), .A2(new_n912), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G952), .B2(G953), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n780), .A2(new_n435), .A3(new_n672), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n848), .B2(KEYINPUT49), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(KEYINPUT49), .B2(new_n848), .ZN(new_n926));
  INV_X1    g740(.A(new_n733), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n718), .A2(new_n926), .A3(new_n927), .A4(new_n815), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n928), .ZN(G75));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n290), .A2(new_n292), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n294), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n934), .A2(new_n938), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n223), .A2(G952), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(G51));
  NAND2_X1  g756(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n921), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n931), .A2(new_n945), .A3(KEYINPUT54), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n622), .B(KEYINPUT57), .Z(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT123), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(new_n950), .A3(new_n946), .A4(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n739), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n932), .A2(new_n803), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n941), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  INV_X1    g769(.A(new_n364), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n941), .ZN(G60));
  INV_X1    g773(.A(new_n941), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n912), .B2(new_n921), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(new_n648), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n944), .A2(new_n946), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n647), .B2(new_n639), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT125), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n931), .A2(new_n688), .A3(new_n686), .A4(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n931), .A2(new_n970), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n960), .B(new_n971), .C1(new_n972), .C2(new_n585), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g790(.A(new_n223), .B1(new_n377), .B2(G224), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n900), .A2(new_n899), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n902), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n980), .B2(new_n223), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n935), .B1(G898), .B2(new_n223), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n981), .B(new_n982), .Z(G69));
  AND4_X1   g797(.A1(new_n792), .A2(new_n897), .A3(new_n721), .A4(new_n783), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n984), .B(new_n829), .C1(new_n821), .C2(new_n822), .ZN(new_n985));
  INV_X1    g799(.A(new_n774), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n986), .B(new_n737), .C1(new_n715), .C2(new_n707), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n734), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n985), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n223), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n490), .B(new_n360), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n810), .A2(new_n721), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n789), .A2(new_n725), .A3(new_n660), .A4(new_n761), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n798), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n829), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n907), .A3(new_n987), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n223), .B1(new_n1000), .B2(new_n823), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n700), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n993), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n995), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1005), .B1(new_n995), .B2(new_n1003), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1006), .A2(new_n1007), .ZN(G72));
  NOR2_X1   g822(.A1(new_n507), .A2(new_n526), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n500), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1000), .A2(new_n823), .A3(new_n980), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OR3_X1    g828(.A1(new_n1011), .A2(KEYINPUT127), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(KEYINPUT127), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1013), .B1(new_n991), .B2(new_n980), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1009), .A2(new_n500), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n508), .A2(new_n527), .A3(new_n509), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n911), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n960), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1017), .A2(new_n1023), .ZN(G57));
endmodule


