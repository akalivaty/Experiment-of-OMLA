//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT17), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n211), .B(KEYINPUT88), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT86), .B(G50gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT85), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G43gat), .B2(G50gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n222), .B2(new_n223), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n218), .B(new_n219), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n212), .B1(new_n214), .B2(KEYINPUT87), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT87), .B2(new_n214), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n209), .B1(new_n210), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n210), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(new_n209), .B2(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT90), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n233), .B(KEYINPUT13), .Z(new_n238));
  OR2_X1    g037(.A1(new_n209), .A2(new_n229), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT91), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n229), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(KEYINPUT91), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT92), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(new_n235), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT11), .B(G169gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT12), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n245), .A3(new_n254), .A4(new_n246), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258));
  XOR2_X1   g057(.A(G15gat), .B(G43gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT67), .ZN(new_n260));
  XNOR2_X1  g059(.A(G71gat), .B(G99gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G227gat), .ZN(new_n263));
  INV_X1    g062(.A(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G169gat), .ZN(new_n266));
  INV_X1    g065(.A(G176gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT65), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(G169gat), .A3(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n266), .A3(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n268), .A2(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n278), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT25), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G183gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT27), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  AND4_X1   g091(.A1(KEYINPUT28), .A2(new_n289), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT27), .B(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n268), .A2(new_n270), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n285), .A2(new_n287), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(G134gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G127gat), .ZN(new_n315));
  INV_X1    g114(.A(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G134gat), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n312), .A2(new_n313), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n317), .ZN(new_n319));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT1), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n303), .A3(new_n302), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT28), .B1(new_n295), .B2(new_n292), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n276), .C1(new_n325), .C2(new_n293), .ZN(new_n326));
  INV_X1    g125(.A(new_n287), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n274), .B2(new_n282), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n326), .B(new_n322), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n265), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n262), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(KEYINPUT66), .A3(KEYINPUT32), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  INV_X1    g134(.A(new_n265), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n321), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n339), .B2(new_n329), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT32), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n331), .B(KEYINPUT32), .C1(new_n332), .C2(new_n262), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n336), .A3(new_n329), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT34), .Z(new_n346));
  AND3_X1   g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n343), .B2(new_n344), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G8gat), .B(G36gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT70), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  INV_X1    g153(.A(G218gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT68), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G197gat), .ZN(new_n363));
  INV_X1    g162(.A(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n357), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(new_n368), .A3(new_n361), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G226gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n264), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n337), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n337), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT69), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI22_X1  g179(.A1(new_n307), .A2(KEYINPUT29), .B1(new_n374), .B2(new_n264), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n373), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n377), .A2(new_n379), .A3(new_n372), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n353), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n381), .B2(new_n376), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n379), .A2(KEYINPUT69), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n372), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n353), .ZN(new_n390));
  INV_X1    g189(.A(new_n385), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n392), .A3(KEYINPUT30), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n384), .A2(new_n385), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n390), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(G22gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n370), .A2(new_n378), .A3(new_n371), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n370), .A2(new_n403), .A3(new_n378), .A4(new_n371), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406));
  INV_X1    g205(.A(G155gat), .ZN(new_n407));
  INV_X1    g206(.A(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(new_n409), .B2(KEYINPUT2), .ZN(new_n410));
  AND2_X1   g209(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n412));
  INV_X1    g211(.A(G141gat), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(G148gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n406), .A2(new_n418), .A3(KEYINPUT2), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G141gat), .B(G148gat), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n418), .B1(new_n406), .B2(KEYINPUT2), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n406), .A2(KEYINPUT71), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(G155gat), .A3(G162gat), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n424), .A2(new_n426), .B1(new_n407), .B2(new_n408), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n417), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n406), .A2(KEYINPUT2), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT72), .ZN(new_n432));
  INV_X1    g231(.A(G148gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G141gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n419), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n427), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n402), .A3(new_n417), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n378), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n372), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT80), .ZN(new_n441));
  INV_X1    g240(.A(G228gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n264), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n444), .A3(new_n372), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n430), .A2(new_n441), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n440), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n433), .ZN(new_n453));
  NAND2_X1  g252(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(G141gat), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n415), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n436), .A2(new_n427), .B1(new_n456), .B2(new_n410), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n400), .B2(new_n402), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n451), .A2(new_n458), .B1(new_n442), .B2(new_n264), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n446), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n450), .B1(new_n446), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n399), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n449), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n450), .A3(new_n459), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n398), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n349), .A2(new_n397), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT0), .ZN(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G85gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n429), .B2(new_n338), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n338), .B1(new_n457), .B2(new_n402), .ZN(new_n476));
  INV_X1    g275(.A(new_n438), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(KEYINPUT76), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n429), .A2(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n438), .A3(new_n338), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(new_n481), .A3(new_n474), .A4(new_n475), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n486), .B2(KEYINPUT5), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n472), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n429), .A2(new_n338), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n457), .A2(new_n322), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n481), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT5), .B1(new_n492), .B2(KEYINPUT74), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n494), .B(new_n481), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  INV_X1    g296(.A(new_n481), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n429), .A2(new_n338), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n437), .A2(new_n417), .B1(new_n318), .B2(new_n321), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n480), .B1(new_n501), .B2(new_n494), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n492), .A2(KEYINPUT74), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n489), .A3(new_n486), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n488), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT77), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n494), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n486), .A2(new_n510), .A3(KEYINPUT5), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT75), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(new_n504), .B1(new_n487), .B2(new_n482), .ZN(new_n513));
  INV_X1    g312(.A(new_n472), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT78), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n482), .A2(new_n487), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n497), .B2(new_n505), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n472), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT77), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n506), .A2(new_n520), .A3(new_n507), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n509), .A2(new_n515), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n512), .A2(new_n504), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n514), .B1(new_n523), .B2(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n468), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n258), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n525), .ZN(new_n529));
  AOI211_X1 g328(.A(KEYINPUT77), .B(KEYINPUT6), .C1(new_n523), .C2(new_n488), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n520), .B1(new_n506), .B2(new_n507), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n515), .A2(new_n519), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT84), .B(KEYINPUT35), .C1(new_n534), .C2(new_n468), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT82), .B1(new_n513), .B2(new_n514), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(new_n507), .A3(new_n538), .A4(new_n506), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  INV_X1    g339(.A(new_n349), .ZN(new_n541));
  INV_X1    g340(.A(new_n467), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n543), .A3(new_n527), .A4(new_n397), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n535), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n397), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n389), .B2(new_n391), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT83), .B1(new_n549), .B2(new_n390), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n394), .A2(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n549), .A2(KEYINPUT83), .A3(new_n390), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT38), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n373), .B1(new_n387), .B2(new_n388), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n377), .A2(new_n379), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n548), .B1(new_n556), .B2(new_n372), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT38), .B(new_n390), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n558), .A2(new_n551), .B1(new_n390), .B2(new_n394), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n554), .A2(new_n525), .A3(new_n539), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n478), .A2(new_n498), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n490), .A2(new_n491), .A3(new_n481), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT39), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(new_n514), .C1(KEYINPUT39), .C2(new_n561), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT40), .Z(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n397), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n537), .A2(new_n538), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n542), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n349), .B(KEYINPUT36), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n547), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n257), .B1(new_n545), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(G57gat), .A2(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G57gat), .A2(G64gat), .ZN(new_n574));
  AND2_X1   g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(KEYINPUT9), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  NOR2_X1   g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n575), .A2(new_n578), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G99gat), .B(G106gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n582), .B1(new_n593), .B2(KEYINPUT99), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT98), .B1(new_n582), .B2(KEYINPUT99), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n581), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n582), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(new_n581), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G230gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n264), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n601), .A2(KEYINPUT100), .A3(KEYINPUT10), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT100), .B1(new_n601), .B2(KEYINPUT10), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n609), .B2(new_n603), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n604), .B(new_n613), .C1(new_n609), .C2(new_n603), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT101), .B1(new_n615), .B2(new_n616), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G127gat), .B(G155gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT20), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n624), .B(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n209), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT95), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n599), .B1(new_n210), .B2(new_n229), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n231), .ZN(new_n638));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT96), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n599), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n645), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n636), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n621), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n572), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n534), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n397), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n202), .B2(new_n661), .ZN(new_n664));
  MUX2_X1   g463(.A(new_n663), .B(new_n664), .S(KEYINPUT42), .Z(G1325gat));
  OR3_X1    g464(.A1(new_n657), .A2(G15gat), .A3(new_n541), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n570), .B(KEYINPUT103), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n657), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n657), .A2(new_n467), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n545), .A2(new_n571), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n650), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n620), .A2(new_n636), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n257), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n534), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n649), .B1(new_n545), .B2(new_n571), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  INV_X1    g481(.A(G29gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n534), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(G1328gat));
  INV_X1    g485(.A(G36gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n682), .A2(new_n687), .A3(new_n546), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n546), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G36gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n697));
  OAI221_X1 g496(.A(new_n692), .B1(new_n690), .B2(new_n688), .C1(new_n696), .C2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n667), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n682), .A2(new_n700), .A3(new_n349), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n678), .A2(KEYINPUT106), .A3(new_n570), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT106), .B1(new_n678), .B2(new_n570), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(G43gat), .A3(new_n706), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n703), .A2(new_n699), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(G1330gat));
  OAI21_X1  g508(.A(new_n220), .B1(new_n678), .B2(new_n467), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n676), .A2(new_n220), .A3(new_n467), .A4(new_n649), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n572), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(KEYINPUT48), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(KEYINPUT107), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT48), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT108), .B(KEYINPUT48), .C1(new_n710), .C2(new_n714), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(G1331gat));
  NOR3_X1   g518(.A1(new_n652), .A2(new_n620), .A3(new_n256), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n673), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n534), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n397), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  NOR3_X1   g528(.A1(new_n721), .A2(G71gat), .A3(new_n541), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n722), .A2(new_n701), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(G71gat), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g532(.A1(new_n721), .A2(new_n467), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(G78gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n673), .A2(KEYINPUT110), .A3(new_n650), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n257), .A2(new_n636), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n681), .A2(KEYINPUT110), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n681), .A2(KEYINPUT110), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n739), .B1(new_n681), .B2(KEYINPUT110), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT111), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n588), .A3(new_n534), .A4(new_n621), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n739), .A2(new_n620), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n675), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n679), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n751), .B2(new_n397), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n620), .A2(G92gat), .A3(new_n397), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n746), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(new_n737), .C1(new_n741), .C2(new_n742), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n762), .A3(new_n756), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n754), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(KEYINPUT52), .ZN(new_n765));
  AOI211_X1 g564(.A(KEYINPUT113), .B(new_n755), .C1(new_n763), .C2(new_n754), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n758), .B1(new_n765), .B2(new_n766), .ZN(G1337gat));
  XOR2_X1   g566(.A(KEYINPUT114), .B(G99gat), .Z(new_n768));
  NOR3_X1   g567(.A1(new_n620), .A2(new_n541), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n751), .B2(new_n667), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1338gat));
  NOR3_X1   g571(.A1(new_n620), .A2(G106gat), .A3(new_n467), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n760), .A2(new_n762), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n775), .A2(new_n542), .A3(new_n776), .A4(new_n750), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n747), .A2(new_n773), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n783), .A3(new_n778), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n774), .B2(new_n778), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n782), .A2(new_n783), .A3(new_n778), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1339gat));
  NOR2_X1   g588(.A1(new_n679), .A2(new_n546), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  INV_X1    g590(.A(new_n636), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n609), .A2(new_n603), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n613), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n609), .A2(new_n603), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT54), .B1(new_n609), .B2(new_n603), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n795), .B(KEYINPUT55), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n242), .A2(new_n238), .A3(new_n243), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n232), .A2(new_n233), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n251), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n255), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(new_n801), .A3(new_n616), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n792), .B1(new_n806), .B2(new_n650), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n618), .B2(new_n619), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n800), .A2(new_n256), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n801), .A2(new_n616), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n808), .B(new_n649), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n620), .A2(new_n257), .A3(new_n651), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n791), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT116), .B(new_n813), .C1(new_n807), .C2(new_n811), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n543), .B(new_n790), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n256), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n814), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n812), .A2(new_n791), .A3(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n543), .A4(new_n790), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n257), .A2(new_n310), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n827), .B2(new_n828), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n308), .A3(new_n621), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n621), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT118), .B1(new_n831), .B2(G120gat), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n833), .B(new_n308), .C1(new_n827), .C2(new_n621), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n830), .B1(new_n832), .B2(new_n834), .ZN(G1341gat));
  OAI21_X1  g634(.A(new_n316), .B1(new_n817), .B2(new_n636), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n792), .A2(G127gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n824), .B2(new_n826), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(G1342gat));
  NOR3_X1   g640(.A1(new_n468), .A2(new_n649), .A3(G134gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n534), .A3(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT56), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n650), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT120), .B1(new_n845), .B2(G134gat), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n847), .B(new_n314), .C1(new_n827), .C2(new_n650), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n667), .A2(new_n542), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n397), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n823), .A2(new_n534), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n413), .A3(new_n256), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n790), .A2(new_n570), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n820), .A2(new_n542), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n542), .C1(new_n815), .C2(new_n816), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n257), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n856), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n411), .A2(new_n412), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n855), .A2(new_n869), .A3(new_n621), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n862), .A2(new_n620), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(KEYINPUT59), .A3(new_n869), .ZN(new_n872));
  XOR2_X1   g671(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n873));
  OAI211_X1 g672(.A(KEYINPUT57), .B(new_n542), .C1(new_n815), .C2(new_n816), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n860), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n857), .A2(new_n620), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n873), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n870), .B1(new_n872), .B2(new_n879), .ZN(G1345gat));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n407), .A3(new_n636), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n854), .A2(new_n636), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT123), .ZN(new_n883));
  AOI21_X1  g682(.A(G155gat), .B1(new_n882), .B2(KEYINPUT123), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n408), .A3(new_n650), .ZN(new_n886));
  OAI21_X1  g685(.A(G162gat), .B1(new_n862), .B2(new_n649), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n534), .A2(new_n397), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n823), .A2(new_n543), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(G169gat), .A3(new_n257), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n890), .B2(new_n257), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n890), .A2(new_n620), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(new_n267), .ZN(G1349gat));
  OAI21_X1  g697(.A(new_n288), .B1(new_n890), .B2(new_n636), .ZN(new_n899));
  INV_X1    g698(.A(new_n543), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n821), .B2(new_n822), .ZN(new_n901));
  INV_X1    g700(.A(new_n295), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n792), .A4(new_n889), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(G1350gat));
  OAI22_X1  g707(.A1(new_n890), .A2(new_n649), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n667), .A2(new_n542), .A3(new_n546), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n679), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n823), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n256), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n667), .A2(new_n889), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n874), .B2(new_n875), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n257), .A2(new_n363), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(new_n920), .ZN(new_n923));
  OAI21_X1  g722(.A(G204gat), .B1(new_n923), .B2(new_n620), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n621), .A2(new_n364), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT62), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n916), .A2(KEYINPUT62), .A3(new_n925), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n354), .A3(new_n792), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n354), .B1(new_n920), .B2(new_n792), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT63), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n923), .B2(new_n649), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n355), .A3(new_n650), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


