

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  INV_X1 U322 ( .A(KEYINPUT115), .ZN(n383) );
  XNOR2_X1 U323 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U324 ( .A(n386), .B(n385), .ZN(n387) );
  NOR2_X1 U325 ( .A1(n409), .A2(n571), .ZN(n410) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n430) );
  XNOR2_X1 U327 ( .A(n431), .B(n430), .ZN(n454) );
  NOR2_X1 U328 ( .A1(n538), .A2(n456), .ZN(n572) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U330 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G176GAT), .B(G183GAT), .Z(n291) );
  XNOR2_X1 U332 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n293) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n295), .B(n294), .Z(n427) );
  XOR2_X1 U338 ( .A(G43GAT), .B(G134GAT), .Z(n404) );
  XOR2_X1 U339 ( .A(G15GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U340 ( .A(n404), .B(n342), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT87), .B(KEYINPUT65), .Z(n297) );
  XNOR2_X1 U342 ( .A(G99GAT), .B(G71GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U345 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n301) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U352 ( .A(G113GAT), .B(n306), .Z(n451) );
  XNOR2_X1 U353 ( .A(n451), .B(KEYINPUT90), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(n427), .B(n309), .Z(n528) );
  INV_X1 U356 ( .A(n528), .ZN(n538) );
  XOR2_X1 U357 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n311) );
  XNOR2_X1 U358 ( .A(G211GAT), .B(KEYINPUT93), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n325) );
  XOR2_X1 U360 ( .A(KEYINPUT22), .B(G218GAT), .Z(n313) );
  XOR2_X1 U361 ( .A(G22GAT), .B(G155GAT), .Z(n334) );
  XOR2_X1 U362 ( .A(G197GAT), .B(KEYINPUT21), .Z(n420) );
  XNOR2_X1 U363 ( .A(n334), .B(n420), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n403) );
  XOR2_X1 U366 ( .A(n314), .B(n403), .Z(n323) );
  XOR2_X1 U367 ( .A(G148GAT), .B(G106GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(G204GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(KEYINPUT74), .B(n317), .Z(n379) );
  XNOR2_X1 U371 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n318), .B(KEYINPUT2), .ZN(n438) );
  XOR2_X1 U373 ( .A(KEYINPUT24), .B(n438), .Z(n320) );
  NAND2_X1 U374 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n379), .B(n321), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n468) );
  XOR2_X1 U379 ( .A(KEYINPUT14), .B(G64GAT), .Z(n327) );
  XNOR2_X1 U380 ( .A(G183GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U382 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U385 ( .A(n331), .B(n330), .Z(n333) );
  XOR2_X1 U386 ( .A(KEYINPUT71), .B(G1GAT), .Z(n348) );
  XOR2_X1 U387 ( .A(G8GAT), .B(G211GAT), .Z(n418) );
  XNOR2_X1 U388 ( .A(n348), .B(n418), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U390 ( .A(n334), .B(KEYINPUT83), .Z(n336) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n338), .B(n337), .Z(n344) );
  XOR2_X1 U394 ( .A(KEYINPUT73), .B(G57GAT), .Z(n340) );
  XNOR2_X1 U395 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U397 ( .A(KEYINPUT72), .B(n341), .Z(n378) );
  XNOR2_X1 U398 ( .A(n342), .B(n378), .ZN(n343) );
  XOR2_X1 U399 ( .A(n344), .B(n343), .Z(n585) );
  XNOR2_X1 U400 ( .A(n585), .B(KEYINPUT114), .ZN(n569) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G197GAT), .Z(n346) );
  XNOR2_X1 U402 ( .A(G36GAT), .B(G22GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n347), .B(G43GAT), .Z(n350) );
  XNOR2_X1 U405 ( .A(n348), .B(G50GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n355) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n351), .B(KEYINPUT7), .ZN(n391) );
  XOR2_X1 U409 ( .A(n391), .B(KEYINPUT29), .Z(n353) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U412 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G113GAT), .Z(n357) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G15GAT), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n359) );
  XNOR2_X1 U417 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n555) );
  INV_X1 U421 ( .A(n555), .ZN(n578) );
  XNOR2_X1 U422 ( .A(G99GAT), .B(G85GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n364), .B(KEYINPUT75), .ZN(n401) );
  XNOR2_X1 U424 ( .A(n401), .B(KEYINPUT33), .ZN(n366) );
  AND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n365) );
  XOR2_X1 U426 ( .A(n366), .B(n365), .Z(n377) );
  XOR2_X1 U427 ( .A(G92GAT), .B(G64GAT), .Z(n417) );
  INV_X1 U428 ( .A(KEYINPUT31), .ZN(n367) );
  NAND2_X1 U429 ( .A1(KEYINPUT76), .A2(n367), .ZN(n370) );
  INV_X1 U430 ( .A(KEYINPUT76), .ZN(n368) );
  NAND2_X1 U431 ( .A1(n368), .A2(KEYINPUT31), .ZN(n369) );
  NAND2_X1 U432 ( .A1(n370), .A2(n369), .ZN(n372) );
  XNOR2_X1 U433 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U435 ( .A(n417), .B(n373), .Z(n375) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(G120GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n581) );
  XOR2_X1 U441 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n382) );
  XOR2_X1 U442 ( .A(n581), .B(n382), .Z(n560) );
  INV_X1 U443 ( .A(n560), .ZN(n541) );
  NAND2_X1 U444 ( .A1(n578), .A2(n541), .ZN(n386) );
  XOR2_X1 U445 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n384) );
  NOR2_X1 U446 ( .A1(n569), .A2(n387), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n388), .B(KEYINPUT117), .ZN(n409) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n390) );
  XNOR2_X1 U449 ( .A(G190GAT), .B(KEYINPUT11), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT9), .B(n391), .Z(n393) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n408) );
  XOR2_X1 U455 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U458 ( .A(n398), .B(G92GAT), .Z(n400) );
  XOR2_X1 U459 ( .A(G36GAT), .B(G218GAT), .Z(n419) );
  XNOR2_X1 U460 ( .A(G106GAT), .B(n419), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n566) );
  INV_X1 U466 ( .A(n566), .ZN(n571) );
  XNOR2_X1 U467 ( .A(n410), .B(KEYINPUT47), .ZN(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT36), .B(n571), .Z(n491) );
  INV_X1 U469 ( .A(n585), .ZN(n563) );
  NOR2_X1 U470 ( .A1(n491), .A2(n563), .ZN(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT45), .B(n411), .ZN(n413) );
  NOR2_X1 U472 ( .A1(n578), .A2(n581), .ZN(n412) );
  NAND2_X1 U473 ( .A1(n413), .A2(n412), .ZN(n414) );
  NAND2_X1 U474 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n416), .B(KEYINPUT48), .ZN(n554) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U479 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n424) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n429) );
  XNOR2_X1 U483 ( .A(n427), .B(G204GAT), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n514) );
  INV_X1 U485 ( .A(n514), .ZN(n526) );
  NAND2_X1 U486 ( .A1(n554), .A2(n526), .ZN(n431) );
  XOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U490 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n435) );
  XNOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT97), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U494 ( .A(G162GAT), .B(n438), .Z(n440) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U499 ( .A(KEYINPUT81), .B(G85GAT), .Z(n445) );
  XNOR2_X1 U500 ( .A(G134GAT), .B(G155GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U503 ( .A(G57GAT), .B(G148GAT), .Z(n449) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(G127GAT), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U507 ( .A(n453), .B(n452), .Z(n524) );
  INV_X1 U508 ( .A(n524), .ZN(n510) );
  NAND2_X1 U509 ( .A1(n454), .A2(n510), .ZN(n462) );
  NOR2_X1 U510 ( .A1(n468), .A2(n462), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n572), .A2(n541), .ZN(n460) );
  XOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XNOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n468), .A2(n538), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT26), .ZN(n552) );
  NOR2_X1 U517 ( .A1(n552), .A2(n462), .ZN(n586) );
  INV_X1 U518 ( .A(n586), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n491), .A2(n463), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT62), .B(n464), .ZN(n465) );
  XOR2_X1 U521 ( .A(G218GAT), .B(n465), .Z(G1355GAT) );
  XOR2_X1 U522 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n483) );
  XOR2_X1 U523 ( .A(KEYINPUT28), .B(n468), .Z(n518) );
  INV_X1 U524 ( .A(n518), .ZN(n530) );
  XNOR2_X1 U525 ( .A(n514), .B(KEYINPUT27), .ZN(n471) );
  OR2_X1 U526 ( .A1(n510), .A2(n471), .ZN(n551) );
  NOR2_X1 U527 ( .A1(n530), .A2(n551), .ZN(n536) );
  XNOR2_X1 U528 ( .A(KEYINPUT91), .B(n528), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n536), .A2(n466), .ZN(n477) );
  NOR2_X1 U530 ( .A1(n538), .A2(n514), .ZN(n467) );
  NOR2_X1 U531 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U532 ( .A(n469), .B(KEYINPUT100), .Z(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(n470), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n552), .A2(n471), .ZN(n472) );
  NOR2_X1 U535 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U536 ( .A(KEYINPUT101), .B(n474), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n475), .A2(n510), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n492) );
  NAND2_X1 U539 ( .A1(n566), .A2(n585), .ZN(n478) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  AND2_X1 U541 ( .A1(n492), .A2(n479), .ZN(n509) );
  NOR2_X1 U542 ( .A1(n555), .A2(n581), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n480), .B(KEYINPUT78), .ZN(n495) );
  NAND2_X1 U544 ( .A1(n509), .A2(n495), .ZN(n481) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(n481), .Z(n488) );
  NAND2_X1 U546 ( .A1(n488), .A2(n524), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n488), .A2(n526), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U552 ( .A1(n528), .A2(n488), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n488), .A2(n530), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n489), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  NOR2_X1 U557 ( .A1(n491), .A2(n585), .ZN(n493) );
  NAND2_X1 U558 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n494), .ZN(n521) );
  NAND2_X1 U560 ( .A1(n495), .A2(n521), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(KEYINPUT106), .ZN(n497) );
  XNOR2_X1 U562 ( .A(KEYINPUT38), .B(n497), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n510), .A2(n505), .ZN(n500) );
  XOR2_X1 U564 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n498), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n514), .A2(n505), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U570 ( .A1(n538), .A2(n505), .ZN(n503) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n518), .A2(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  NOR2_X1 U577 ( .A1(n578), .A2(n560), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(n509), .ZN(n517) );
  NOR2_X1 U579 ( .A1(n510), .A2(n517), .ZN(n512) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NOR2_X1 U583 ( .A1(n514), .A2(n517), .ZN(n515) );
  XOR2_X1 U584 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U585 ( .A1(n538), .A2(n517), .ZN(n516) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT111), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n526), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n528), .A2(n531), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n533) );
  NAND2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n554), .A2(n536), .ZN(n537) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n548), .A2(n578), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(KEYINPUT118), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n543) );
  NAND2_X1 U609 ( .A1(n548), .A2(n541), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n569), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n571), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n565) );
  NOR2_X1 U621 ( .A1(n555), .A2(n565), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n565), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n578), .A2(n572), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n574), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(n577), .Z(n580) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n586), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
endmodule

