

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(G2104), .A2(n523), .ZN(n886) );
  NOR2_X1 U557 ( .A1(n948), .A2(n610), .ZN(n609) );
  NOR2_X1 U558 ( .A1(n533), .A2(n532), .ZN(G160) );
  OR2_X1 U559 ( .A1(n707), .A2(n706), .ZN(n520) );
  NAND2_X1 U560 ( .A1(n700), .A2(n699), .ZN(n521) );
  INV_X1 U561 ( .A(KEYINPUT28), .ZN(n608) );
  AND2_X1 U562 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U563 ( .A1(n711), .A2(n602), .ZN(n674) );
  NAND2_X1 U564 ( .A1(G160), .A2(G40), .ZN(n710) );
  AND2_X1 U565 ( .A1(n708), .A2(n520), .ZN(n709) );
  NOR2_X1 U566 ( .A1(G651), .A2(n551), .ZN(n794) );
  INV_X1 U567 ( .A(G2105), .ZN(n523) );
  AND2_X1 U568 ( .A1(n523), .A2(G2104), .ZN(n879) );
  NAND2_X1 U569 ( .A1(G101), .A2(n879), .ZN(n522) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n522), .Z(n526) );
  NAND2_X1 U571 ( .A1(G125), .A2(n886), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT65), .B(n524), .Z(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n533) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U575 ( .A1(G113), .A2(n884), .ZN(n531) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X2 U579 ( .A(KEYINPUT66), .B(n529), .ZN(n880) );
  NAND2_X1 U580 ( .A1(G137), .A2(n880), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U582 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n535) );
  XOR2_X1 U583 ( .A(G651), .B(KEYINPUT68), .Z(n550) );
  NOR2_X1 U584 ( .A1(G543), .A2(n550), .ZN(n534) );
  XNOR2_X1 U585 ( .A(n535), .B(n534), .ZN(n793) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n551) );
  NAND2_X1 U587 ( .A1(G87), .A2(n551), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G74), .A2(G651), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n793), .A2(n538), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G49), .A2(n794), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT85), .B(n539), .Z(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(G288) );
  AND2_X1 U594 ( .A1(n880), .A2(G138), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n879), .A2(G102), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G114), .A2(n884), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT91), .B(n542), .Z(n543) );
  AND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n886), .A2(G126), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G53), .A2(n794), .ZN(n549) );
  XNOR2_X1 U603 ( .A(n549), .B(KEYINPUT72), .ZN(n559) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n789) );
  NAND2_X1 U605 ( .A1(G78), .A2(n789), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G65), .A2(n793), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n557) );
  NOR2_X1 U608 ( .A1(G543), .A2(G651), .ZN(n554) );
  XNOR2_X1 U609 ( .A(n554), .B(KEYINPUT64), .ZN(n790) );
  NAND2_X1 U610 ( .A1(G91), .A2(n790), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT71), .B(n555), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U614 ( .A1(G64), .A2(n793), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G52), .A2(n794), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n789), .A2(G77), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G90), .A2(n790), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U621 ( .A1(n566), .A2(n565), .ZN(G171) );
  INV_X1 U622 ( .A(G171), .ZN(G301) );
  NAND2_X1 U623 ( .A1(n789), .A2(G76), .ZN(n567) );
  XNOR2_X1 U624 ( .A(KEYINPUT78), .B(n567), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G89), .A2(n790), .ZN(n568) );
  XNOR2_X1 U626 ( .A(KEYINPUT4), .B(n568), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n571), .B(KEYINPUT5), .ZN(n576) );
  NAND2_X1 U629 ( .A1(G63), .A2(n793), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G51), .A2(n794), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U634 ( .A(n577), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .ZN(n578) );
  XNOR2_X1 U636 ( .A(n578), .B(KEYINPUT79), .ZN(G286) );
  NAND2_X1 U637 ( .A1(n789), .A2(G75), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G88), .A2(n790), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U640 ( .A(KEYINPUT89), .B(n581), .ZN(n587) );
  NAND2_X1 U641 ( .A1(G62), .A2(n793), .ZN(n582) );
  XNOR2_X1 U642 ( .A(n582), .B(KEYINPUT87), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G50), .A2(n794), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT88), .B(n583), .Z(n584) );
  NOR2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G303) );
  INV_X1 U647 ( .A(G303), .ZN(G166) );
  NAND2_X1 U648 ( .A1(G61), .A2(n793), .ZN(n588) );
  XNOR2_X1 U649 ( .A(n588), .B(KEYINPUT86), .ZN(n595) );
  NAND2_X1 U650 ( .A1(n794), .A2(G48), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G86), .A2(n790), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U653 ( .A1(n789), .A2(G73), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT2), .B(n591), .Z(n592) );
  NOR2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(G305) );
  NAND2_X1 U657 ( .A1(n793), .A2(G60), .ZN(n597) );
  NAND2_X1 U658 ( .A1(G85), .A2(n790), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G72), .A2(n789), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G47), .A2(n794), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n600) );
  OR2_X1 U663 ( .A1(n601), .A2(n600), .ZN(G290) );
  AND2_X1 U664 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NOR2_X1 U665 ( .A1(G1976), .A2(G288), .ZN(n947) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n711) );
  INV_X1 U667 ( .A(n710), .ZN(n602) );
  NOR2_X1 U668 ( .A1(G2084), .A2(n674), .ZN(n657) );
  NAND2_X1 U669 ( .A1(G8), .A2(n657), .ZN(n672) );
  NAND2_X1 U670 ( .A1(G8), .A2(n674), .ZN(n707) );
  NOR2_X1 U671 ( .A1(G1966), .A2(n707), .ZN(n670) );
  INV_X1 U672 ( .A(G299), .ZN(n948) );
  XOR2_X1 U673 ( .A(KEYINPUT98), .B(n674), .Z(n636) );
  NAND2_X1 U674 ( .A1(G2072), .A2(n636), .ZN(n604) );
  INV_X1 U675 ( .A(KEYINPUT27), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U677 ( .A(n636), .ZN(n650) );
  NAND2_X1 U678 ( .A1(G1956), .A2(n650), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT101), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n609), .B(n608), .ZN(n646) );
  NAND2_X1 U682 ( .A1(n948), .A2(n610), .ZN(n644) );
  NAND2_X1 U683 ( .A1(n793), .A2(G66), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n611), .Z(n613) );
  NAND2_X1 U685 ( .A1(G92), .A2(n790), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G79), .A2(n789), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G54), .A2(n794), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U692 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(n946) );
  NAND2_X1 U694 ( .A1(n793), .A2(G56), .ZN(n621) );
  XOR2_X1 U695 ( .A(KEYINPUT14), .B(n621), .Z(n627) );
  NAND2_X1 U696 ( .A1(G81), .A2(n790), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT12), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G68), .A2(n789), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U700 ( .A(KEYINPUT13), .B(n625), .Z(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n628), .B(KEYINPUT74), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G43), .A2(n794), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n961) );
  INV_X1 U705 ( .A(n674), .ZN(n652) );
  AND2_X1 U706 ( .A1(n652), .A2(G1996), .ZN(n631) );
  XOR2_X1 U707 ( .A(n631), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U708 ( .A1(n674), .A2(G1341), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n961), .A2(n634), .ZN(n635) );
  OR2_X1 U711 ( .A1(n946), .A2(n635), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n946), .A2(n635), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G2067), .A2(n636), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G1348), .A2(n674), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n656) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT99), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT25), .ZN(n1000) );
  NOR2_X1 U724 ( .A1(n1000), .A2(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT100), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n652), .A2(G1961), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n663) );
  OR2_X1 U728 ( .A1(n663), .A2(G301), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n668) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n660) );
  NOR2_X1 U731 ( .A1(n670), .A2(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n658), .A2(G8), .ZN(n659) );
  XOR2_X1 U733 ( .A(n660), .B(n659), .Z(n661) );
  NOR2_X1 U734 ( .A1(G168), .A2(n661), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT104), .B(n662), .Z(n665) );
  NAND2_X1 U736 ( .A1(n663), .A2(G301), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT31), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n673) );
  INV_X1 U740 ( .A(n673), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n673), .A2(G286), .ZN(n681) );
  INV_X1 U744 ( .A(G8), .ZN(n679) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n707), .ZN(n676) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n674), .ZN(n675) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U748 ( .A1(n677), .A2(G303), .ZN(n678) );
  OR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT32), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n703) );
  INV_X1 U752 ( .A(G1971), .ZN(n979) );
  NAND2_X1 U753 ( .A1(G166), .A2(n979), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n703), .A2(n685), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n947), .A2(n686), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n952), .A2(n687), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n694), .A2(KEYINPUT105), .ZN(n690) );
  NAND2_X1 U758 ( .A1(KEYINPUT33), .A2(n947), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT106), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  INV_X1 U761 ( .A(n707), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n691), .A2(n693), .ZN(n700) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n943) );
  NAND2_X1 U764 ( .A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(n692) );
  AND2_X1 U765 ( .A1(n943), .A2(n692), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n696) );
  NOR2_X1 U767 ( .A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U771 ( .A1(G8), .A2(n701), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n704), .A2(n707), .ZN(n708) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XOR2_X1 U775 ( .A(n705), .B(KEYINPUT24), .Z(n706) );
  NAND2_X1 U776 ( .A1(n521), .A2(n709), .ZN(n746) );
  XNOR2_X1 U777 ( .A(G1986), .B(G290), .ZN(n951) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n758) );
  NAND2_X1 U779 ( .A1(n951), .A2(n758), .ZN(n712) );
  XNOR2_X1 U780 ( .A(n712), .B(KEYINPUT92), .ZN(n725) );
  NAND2_X1 U781 ( .A1(G104), .A2(n879), .ZN(n714) );
  NAND2_X1 U782 ( .A1(G140), .A2(n880), .ZN(n713) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n715), .ZN(n721) );
  NAND2_X1 U785 ( .A1(n884), .A2(G116), .ZN(n716) );
  XOR2_X1 U786 ( .A(KEYINPUT93), .B(n716), .Z(n718) );
  NAND2_X1 U787 ( .A1(n886), .A2(G128), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U789 ( .A(n719), .B(KEYINPUT35), .Z(n720) );
  NOR2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U791 ( .A(KEYINPUT36), .B(n722), .Z(n723) );
  XOR2_X1 U792 ( .A(KEYINPUT94), .B(n723), .Z(n892) );
  XNOR2_X1 U793 ( .A(KEYINPUT37), .B(G2067), .ZN(n756) );
  OR2_X1 U794 ( .A1(n892), .A2(n756), .ZN(n724) );
  XNOR2_X1 U795 ( .A(n724), .B(KEYINPUT95), .ZN(n924) );
  NAND2_X1 U796 ( .A1(n758), .A2(n924), .ZN(n754) );
  NAND2_X1 U797 ( .A1(n725), .A2(n754), .ZN(n744) );
  NAND2_X1 U798 ( .A1(G107), .A2(n884), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G95), .A2(n879), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U801 ( .A1(n886), .A2(G119), .ZN(n728) );
  XOR2_X1 U802 ( .A(KEYINPUT96), .B(n728), .Z(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G131), .A2(n880), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n869) );
  NAND2_X1 U806 ( .A1(G1991), .A2(n869), .ZN(n741) );
  NAND2_X1 U807 ( .A1(G117), .A2(n884), .ZN(n734) );
  NAND2_X1 U808 ( .A1(G129), .A2(n886), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n879), .A2(G105), .ZN(n735) );
  XOR2_X1 U811 ( .A(KEYINPUT38), .B(n735), .Z(n736) );
  NOR2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U813 ( .A1(G141), .A2(n880), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n863) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n863), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n925) );
  NAND2_X1 U817 ( .A1(n758), .A2(n925), .ZN(n742) );
  XNOR2_X1 U818 ( .A(KEYINPUT97), .B(n742), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n761) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n863), .ZN(n747) );
  XOR2_X1 U822 ( .A(KEYINPUT107), .B(n747), .Z(n928) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n869), .ZN(n748) );
  XOR2_X1 U824 ( .A(KEYINPUT109), .B(n748), .Z(n934) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n749) );
  XNOR2_X1 U826 ( .A(KEYINPUT108), .B(n749), .ZN(n750) );
  NOR2_X1 U827 ( .A1(n934), .A2(n750), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n751), .A2(n925), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n928), .A2(n752), .ZN(n753) );
  XNOR2_X1 U830 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U832 ( .A1(n892), .A2(n756), .ZN(n921) );
  NAND2_X1 U833 ( .A1(n757), .A2(n921), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  NAND2_X1 U840 ( .A1(G94), .A2(G452), .ZN(n763) );
  XOR2_X1 U841 ( .A(KEYINPUT70), .B(n763), .Z(G173) );
  XOR2_X1 U842 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n765) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U844 ( .A(n765), .B(n764), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n822) );
  NAND2_X1 U846 ( .A1(n822), .A2(G567), .ZN(n766) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U848 ( .A(G860), .ZN(n829) );
  OR2_X1 U849 ( .A1(n961), .A2(n829), .ZN(G153) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n768) );
  OR2_X1 U851 ( .A1(n946), .A2(G868), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n769) );
  XNOR2_X1 U854 ( .A(n769), .B(KEYINPUT80), .ZN(n771) );
  INV_X1 U855 ( .A(G868), .ZN(n807) );
  NOR2_X1 U856 ( .A1(n807), .A2(G286), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n829), .A2(G559), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n772), .A2(n946), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n961), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G868), .A2(n946), .ZN(n774) );
  NOR2_X1 U863 ( .A1(G559), .A2(n774), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT81), .B(n777), .Z(G282) );
  XNOR2_X1 U866 ( .A(G2100), .B(KEYINPUT83), .ZN(n787) );
  NAND2_X1 U867 ( .A1(G123), .A2(n886), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n778), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G111), .A2(n884), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(KEYINPUT82), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G99), .A2(n879), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G135), .A2(n880), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n926) );
  XNOR2_X1 U876 ( .A(n926), .B(G2096), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n946), .ZN(n788) );
  XOR2_X1 U879 ( .A(n961), .B(n788), .Z(n828) );
  NAND2_X1 U880 ( .A1(n789), .A2(G80), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G93), .A2(n790), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT84), .B(n799), .Z(n830) );
  XNOR2_X1 U888 ( .A(G166), .B(n830), .ZN(n805) );
  XNOR2_X1 U889 ( .A(KEYINPUT90), .B(G305), .ZN(n800) );
  XNOR2_X1 U890 ( .A(n800), .B(G288), .ZN(n801) );
  XNOR2_X1 U891 ( .A(KEYINPUT19), .B(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(G290), .B(n948), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n805), .B(n804), .ZN(n896) );
  XNOR2_X1 U895 ( .A(n828), .B(n896), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n806), .A2(G868), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n807), .A2(n830), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n810) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U907 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U908 ( .A1(G96), .A2(n816), .ZN(n826) );
  NAND2_X1 U909 ( .A1(n826), .A2(G2106), .ZN(n820) );
  NAND2_X1 U910 ( .A1(G120), .A2(G69), .ZN(n817) );
  NOR2_X1 U911 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U912 ( .A1(G108), .A2(n818), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n827), .A2(G567), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n832) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n832), .A2(n821), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U920 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G325) );
  XOR2_X1 U925 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(G145) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(n832), .ZN(G319) );
  XNOR2_X1 U932 ( .A(G1996), .B(KEYINPUT41), .ZN(n842) );
  XOR2_X1 U933 ( .A(G1971), .B(G1961), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1986), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U936 ( .A(G1976), .B(G1981), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1966), .B(G1956), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2474), .B(KEYINPUT116), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(G229) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n843), .B(KEYINPUT42), .ZN(n853) );
  XOR2_X1 U945 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2678), .B(G2100), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G2096), .B(G2084), .Z(n847) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2072), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G124), .A2(n886), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n884), .A2(G112), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G100), .A2(n879), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G136), .A2(n880), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT119), .B(KEYINPUT46), .Z(n862) );
  XNOR2_X1 U964 ( .A(n926), .B(KEYINPUT48), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n863), .B(G162), .ZN(n865) );
  XNOR2_X1 U967 ( .A(G164), .B(G160), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G118), .A2(n884), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G130), .A2(n886), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n879), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G142), .A2(n880), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(n878), .B(n877), .Z(n894) );
  NAND2_X1 U980 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(KEYINPUT117), .B(n883), .Z(n891) );
  NAND2_X1 U984 ( .A1(n884), .A2(G115), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(KEYINPUT118), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n917) );
  XNOR2_X1 U990 ( .A(n892), .B(n917), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n961), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(G171), .B(n946), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U996 ( .A(G286), .B(n899), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U998 ( .A(G2443), .B(G2451), .Z(n902) );
  XNOR2_X1 U999 ( .A(G2446), .B(G2454), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n903), .B(G2427), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1004 ( .A(G2435), .B(KEYINPUT110), .Z(n907) );
  XNOR2_X1 U1005 ( .A(G2430), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n909), .B(n908), .Z(n910) );
  NAND2_X1 U1008 ( .A1(G14), .A2(n910), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1018 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1023) );
  INV_X1 U1019 ( .A(KEYINPUT55), .ZN(n941) );
  XOR2_X1 U1020 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(n920), .B(KEYINPUT50), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n937) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G160), .B(G2084), .Z(n931) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT120), .B(n938), .ZN(n939) );
  XOR2_X1 U1036 ( .A(KEYINPUT52), .B(n939), .Z(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .ZN(n967) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G168), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(n945), .B(KEYINPUT57), .ZN(n965) );
  XNOR2_X1 U1043 ( .A(n946), .B(G1348), .ZN(n960) );
  XOR2_X1 U1044 ( .A(n947), .B(KEYINPUT122), .Z(n950) );
  XNOR2_X1 U1045 ( .A(n948), .B(G1956), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n958) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G301), .B(G1961), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G303), .B(G1971), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G1341), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n996) );
  INV_X1 U1058 ( .A(G16), .ZN(n994) );
  XOR2_X1 U1059 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n992) );
  XNOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(G4), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G1956), .B(G20), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1066 ( .A(KEYINPUT123), .B(G1981), .Z(n973) );
  XNOR2_X1 U1067 ( .A(G6), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1070 ( .A(G1961), .B(G5), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n990) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G21), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1976), .B(G23), .ZN(n983) );
  XOR2_X1 U1074 ( .A(G1986), .B(G24), .Z(n981) );
  XNOR2_X1 U1075 ( .A(n979), .B(G22), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(n985), .B(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n992), .B(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1019) );
  XOR2_X1 U1086 ( .A(G1991), .B(G25), .Z(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G2067), .B(G26), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G33), .B(G2072), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1996), .B(G32), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G27), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT53), .B(n1007), .Z(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT54), .B(G34), .Z(n1008) );
  XNOR2_X1 U1098 ( .A(G2084), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G35), .B(G2090), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT55), .B(n1013), .ZN(n1015) );
  INV_X1 U1103 ( .A(G29), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(KEYINPUT121), .B(n1017), .Z(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1023), .B(n1022), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

