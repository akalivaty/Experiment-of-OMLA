//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT77), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT18), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  OR2_X1    g0050(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n208), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n218), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n255), .A2(new_n260), .B1(new_n259), .B2(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT16), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT75), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT7), .B1(new_n269), .B2(new_n209), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n271), .B(G20), .C1(new_n266), .C2(new_n268), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n264), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(G20), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT75), .B1(new_n275), .B2(KEYINPUT7), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n263), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n209), .A2(new_n265), .A3(KEYINPUT67), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G20), .B2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G159), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n250), .A2(new_n263), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n283), .B2(new_n201), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n262), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n267), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n288));
  OAI211_X1 g0088(.A(KEYINPUT7), .B(new_n209), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n275), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(G68), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n258), .B1(new_n291), .B2(KEYINPUT16), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n261), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n266), .A2(new_n268), .A3(G226), .A4(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n266), .A2(new_n268), .A3(G223), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G87), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(G1), .A2(G13), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G41), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n208), .A2(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n304), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n306), .A2(G232), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n300), .A2(G179), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n310), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n305), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(G232), .A3(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n299), .B2(new_n298), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT76), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n312), .B(new_n321), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n248), .B(new_n249), .C1(new_n293), .C2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n249), .B1(new_n293), .B2(new_n323), .ZN(new_n325));
  INV_X1    g0125(.A(new_n261), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT75), .B1(new_n275), .B2(new_n289), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n269), .A2(new_n209), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n264), .B1(new_n328), .B2(new_n271), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n285), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT16), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n270), .B2(new_n272), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n257), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n326), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n336), .A2(KEYINPUT18), .A3(new_n320), .A4(new_n322), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n325), .A2(KEYINPUT77), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT17), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n300), .A2(new_n340), .A3(new_n341), .A4(new_n311), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G200), .B2(new_n317), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n317), .B2(new_n341), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n339), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n286), .A2(new_n292), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n300), .A2(new_n311), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT78), .B1(new_n348), .B2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(G200), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n351), .A3(new_n342), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n347), .A2(KEYINPUT17), .A3(new_n326), .A4(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n346), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT79), .B1(new_n346), .B2(new_n353), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n324), .B(new_n338), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n281), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT66), .B1(new_n265), .B2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT66), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n209), .A3(G33), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n253), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n258), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n254), .A2(G50), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n260), .A2(new_n364), .B1(G50), .B2(new_n259), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n274), .A2(G222), .A3(new_n295), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n274), .A2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G223), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n367), .B1(new_n368), .B2(new_n274), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n299), .ZN(new_n372));
  INV_X1    g0172(.A(new_n313), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G226), .B2(new_n306), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n366), .B1(new_n375), .B2(new_n318), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G179), .B2(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n372), .A2(G190), .A3(new_n374), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT9), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n366), .B(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n382), .A2(new_n379), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n379), .A3(new_n383), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT10), .A3(new_n381), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n378), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n306), .A2(G238), .B1(new_n308), .B2(new_n310), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n274), .A2(G226), .A3(new_n295), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n299), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT13), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n341), .B1(new_n398), .B2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n299), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n392), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT72), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n400), .A2(new_n401), .A3(new_n404), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n209), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n361), .B2(G77), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n281), .A2(G50), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n258), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n402), .A2(new_n399), .A3(new_n392), .ZN(new_n419));
  OAI21_X1  g0219(.A(G200), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(KEYINPUT73), .A3(new_n415), .ZN(new_n421));
  INV_X1    g0221(.A(G13), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(G1), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT12), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n410), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n423), .A2(new_n410), .A3(new_n424), .A4(new_n425), .ZN(new_n428));
  INV_X1    g0228(.A(new_n260), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n263), .B1(new_n208), .B2(G20), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n418), .A2(new_n420), .A3(new_n421), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n409), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G169), .B1(new_n419), .B2(new_n403), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(G179), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n419), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n400), .A3(new_n404), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(G169), .C1(new_n419), .C2(new_n403), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n418), .A2(new_n421), .A3(new_n431), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n434), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n274), .A2(G232), .A3(new_n295), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  INV_X1    g0247(.A(G238), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n446), .B1(new_n447), .B2(new_n274), .C1(new_n369), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n299), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n373), .B1(G244), .B2(new_n306), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G179), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n318), .B2(new_n452), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n361), .B1(G20), .B2(G77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n253), .A2(new_n281), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n258), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g0259(.A(new_n459), .B(KEYINPUT68), .Z(new_n460));
  AOI21_X1  g0260(.A(new_n368), .B1(new_n208), .B2(G20), .ZN(new_n461));
  OR3_X1    g0261(.A1(new_n259), .A2(KEYINPUT69), .A3(G77), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT69), .B1(new_n259), .B2(G77), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n429), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n452), .A2(G200), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n341), .B2(new_n452), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n356), .A2(new_n390), .A3(new_n445), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n266), .A2(new_n268), .A3(new_n209), .A4(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT22), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n274), .A2(new_n473), .A3(new_n209), .A4(G87), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G20), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n209), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n447), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n475), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n476), .B1(new_n475), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n257), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n208), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n259), .A2(new_n486), .A3(new_n218), .A4(new_n256), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n259), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(KEYINPUT25), .A3(new_n447), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT25), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n259), .B2(G107), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n488), .A2(G107), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n266), .A2(new_n268), .A3(G257), .A4(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n266), .A2(new_n268), .A3(G250), .A4(new_n295), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G294), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n314), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT86), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n208), .A2(G45), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n299), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n500), .A2(new_n501), .B1(G264), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n308), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n437), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n498), .A2(new_n499), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n299), .A3(new_n501), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(G264), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n508), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n318), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n494), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(G200), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n511), .A2(G190), .A3(new_n512), .A4(new_n508), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n485), .A3(new_n493), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n506), .A2(G270), .B1(new_n308), .B2(new_n505), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n266), .A2(new_n268), .A3(G264), .A4(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n266), .A2(new_n268), .A3(G257), .A4(new_n295), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n274), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n299), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(G179), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n318), .B1(new_n524), .B2(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n256), .A2(new_n218), .B1(G20), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n209), .C1(G33), .C2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n259), .A2(G116), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n487), .B2(new_n535), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT84), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(new_n539), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n543), .B1(new_n488), .B2(G116), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n534), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n555), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n524), .A2(new_n529), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n559), .C1(new_n341), .C2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n555), .A2(new_n531), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n533), .ZN(new_n563));
  AOI211_X1 g0363(.A(KEYINPUT85), .B(KEYINPUT21), .C1(new_n555), .C2(new_n531), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n556), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n259), .A2(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n488), .B2(G97), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n538), .A2(new_n447), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n205), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n538), .A2(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n209), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n368), .B1(new_n278), .B2(new_n280), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(KEYINPUT80), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(KEYINPUT80), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(G107), .B1(new_n327), .B2(new_n329), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT82), .B(new_n568), .C1(new_n583), .C2(new_n258), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n258), .B1(new_n581), .B2(new_n582), .ZN(new_n586));
  INV_X1    g0386(.A(new_n568), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT5), .B(G41), .ZN(new_n589));
  INV_X1    g0389(.A(new_n502), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G257), .A3(new_n314), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n508), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(new_n295), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n295), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n537), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n593), .B1(new_n299), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n341), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(G200), .B2(new_n600), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n584), .A2(new_n588), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n568), .B1(new_n583), .B2(new_n258), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G179), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n318), .B2(new_n600), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n308), .A2(new_n590), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n314), .A2(G250), .A3(new_n502), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n266), .A2(new_n268), .A3(G238), .A4(new_n295), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n477), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(new_n299), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n350), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(G190), .B2(new_n614), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n274), .A2(new_n209), .A3(G68), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n209), .B1(new_n396), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G87), .B2(new_n206), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT19), .B1(new_n361), .B2(G97), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n257), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n455), .A2(new_n489), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(G87), .B2(new_n488), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n613), .A2(new_n299), .ZN(new_n627));
  INV_X1    g0427(.A(new_n610), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G169), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n437), .B2(new_n629), .ZN(new_n631));
  XOR2_X1   g0431(.A(new_n455), .B(KEYINPUT83), .Z(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n623), .B(new_n624), .C1(new_n633), .C2(new_n487), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n616), .A2(new_n626), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n603), .A2(new_n607), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n470), .A2(new_n523), .A3(new_n566), .A4(new_n636), .ZN(G372));
  XNOR2_X1  g0437(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n336), .A2(new_n319), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n336), .B2(new_n319), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n346), .A2(new_n353), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT79), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n346), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n432), .B1(new_n406), .B2(new_n408), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n444), .B1(new_n647), .B2(new_n466), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(new_n386), .B2(new_n388), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n378), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n603), .A2(new_n607), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n616), .A2(new_n626), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n515), .B(new_n556), .C1(new_n563), .C2(new_n564), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n518), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n631), .A2(new_n660), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n634), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n607), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(KEYINPUT26), .A3(new_n635), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n584), .A2(new_n588), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n663), .A2(new_n606), .A3(new_n667), .A4(new_n657), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n470), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n654), .A2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n423), .A2(new_n209), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT91), .ZN(new_n677));
  INV_X1    g0477(.A(G213), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n675), .B2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n557), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n565), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n556), .B1(new_n563), .B2(new_n564), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n674), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n494), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n523), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n515), .A2(new_n682), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n682), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n521), .B2(new_n522), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n515), .A2(new_n689), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n212), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n216), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n507), .A2(new_n600), .A3(new_n614), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n530), .A2(KEYINPUT92), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n524), .A2(new_n529), .A3(new_n709), .A4(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n710), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n507), .A2(new_n600), .A3(new_n614), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n558), .A2(new_n629), .A3(new_n437), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n600), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n513), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT93), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n689), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n523), .A2(new_n566), .A3(new_n636), .A4(new_n682), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n682), .C1(new_n664), .C2(new_n670), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n665), .A2(new_n669), .A3(new_n635), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n659), .A3(new_n663), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n732), .B1(new_n737), .B2(new_n682), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n706), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n422), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n208), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n701), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n688), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n685), .A2(new_n674), .A3(new_n687), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n685), .A2(new_n687), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n212), .A2(new_n274), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n212), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n274), .B(new_n700), .C1(new_n302), .C2(new_n217), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n243), .A2(G45), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n218), .B1(G20), .B2(new_n318), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n745), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  INV_X1    g0563(.A(new_n759), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n209), .A2(new_n437), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(new_n350), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n209), .A2(G179), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n767), .A2(G322), .B1(new_n771), .B2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(new_n341), .A3(G200), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n772), .B1(new_n773), .B2(new_n774), .C1(new_n778), .C2(new_n527), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n765), .A2(new_n769), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n765), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT33), .B(G317), .Z(new_n785));
  OAI221_X1 g0585(.A(new_n269), .B1(new_n780), .B2(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(new_n341), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n209), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n779), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n796));
  INV_X1    g0596(.A(G87), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n778), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n274), .B1(new_n774), .B2(new_n447), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n766), .A2(new_n250), .B1(new_n780), .B2(new_n368), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G97), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT95), .B(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n770), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT32), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G50), .A2(new_n787), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n808), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(KEYINPUT32), .B1(new_n783), .B2(G68), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n801), .A2(new_n806), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n796), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n752), .B(new_n763), .C1(new_n764), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n748), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n671), .A2(new_n682), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n465), .A2(new_n468), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n682), .B1(new_n460), .B2(new_n464), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n466), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n454), .A2(new_n465), .A3(new_n682), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n824), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n682), .B(new_n826), .C1(new_n664), .C2(new_n670), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n745), .B1(new_n829), .B2(new_n730), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n730), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n780), .ZN(new_n832));
  INV_X1    g0632(.A(new_n807), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n767), .A2(G143), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n784), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G137), .B2(new_n787), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n839));
  INV_X1    g0639(.A(new_n774), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n269), .B1(new_n840), .B2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n250), .B2(new_n792), .C1(new_n842), .C2(new_n770), .ZN(new_n843));
  INV_X1    g0643(.A(new_n778), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(G50), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n269), .B1(new_n770), .B2(new_n781), .C1(new_n788), .C2(new_n527), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G283), .B2(new_n783), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(G107), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n766), .A2(new_n790), .B1(new_n774), .B2(new_n797), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G116), .B2(new_n832), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n806), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n759), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n745), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n759), .A2(new_n749), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n368), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n856), .B(new_n859), .C1(new_n750), .C2(new_n826), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n831), .A2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n742), .A2(new_n208), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n291), .A2(KEYINPUT16), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n261), .B1(new_n863), .B2(new_n292), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n680), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n356), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n320), .A2(new_n322), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n336), .B1(new_n867), .B2(new_n681), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT37), .B1(new_n293), .B2(new_n352), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n681), .A2(new_n319), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n336), .A2(new_n345), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n868), .A2(new_n869), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n875), .B(new_n872), .C1(new_n356), .C2(new_n865), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT39), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n866), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n336), .B2(new_n345), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n336), .B1(new_n319), .B2(new_n681), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n347), .A2(KEYINPUT102), .A3(new_n326), .A4(new_n352), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n868), .A2(new_n869), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n293), .A2(new_n680), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n641), .B2(new_n642), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n878), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n877), .A2(KEYINPUT101), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n444), .A2(new_n689), .ZN(new_n894));
  INV_X1    g0694(.A(new_n865), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n338), .A2(new_n324), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n646), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n875), .B1(new_n897), .B2(new_n872), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n878), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT101), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT39), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n893), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n443), .B(new_n689), .C1(new_n647), .C2(new_n442), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n443), .A2(new_n689), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n434), .A2(new_n444), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n827), .B2(new_n823), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n908), .A2(new_n899), .B1(new_n641), .B2(new_n680), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n470), .B1(new_n734), .B2(new_n738), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n654), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n720), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n727), .A2(new_n914), .A3(new_n725), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n824), .B1(new_n903), .B2(new_n905), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(new_n876), .C2(new_n889), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n917), .A2(KEYINPUT40), .B1(new_n899), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n470), .A2(new_n915), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n674), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(KEYINPUT103), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT103), .B2(new_n923), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n862), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n913), .B2(new_n925), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n573), .A2(new_n576), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT35), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT35), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(G116), .A3(new_n219), .A4(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n216), .A2(new_n368), .A3(new_n283), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(KEYINPUT100), .B1(new_n202), .B2(G68), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(KEYINPUT100), .B2(new_n934), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n422), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(new_n933), .A3(new_n937), .ZN(G367));
  NOR2_X1   g0738(.A1(new_n700), .A2(new_n274), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n238), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n760), .C1(new_n212), .C2(new_n455), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n269), .B1(new_n780), .B2(new_n773), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n788), .A2(new_n781), .B1(new_n447), .B2(new_n792), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(G294), .C2(new_n783), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n766), .A2(new_n527), .B1(new_n774), .B2(new_n538), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G317), .B2(new_n771), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n778), .B2(new_n535), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n844), .A2(KEYINPUT46), .A3(G116), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n944), .A2(new_n946), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n766), .A2(new_n835), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n274), .B1(new_n774), .B2(new_n368), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT107), .B(G137), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n951), .B(new_n952), .C1(new_n771), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(G143), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n250), .B2(new_n778), .C1(new_n955), .C2(new_n788), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n805), .A2(G68), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n783), .A2(new_n833), .B1(new_n832), .B2(G50), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT106), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(KEYINPUT106), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n950), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  OAI211_X1 g0763(.A(new_n745), .B(new_n941), .C1(new_n963), .C2(new_n764), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT108), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n663), .A2(new_n657), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n682), .A2(new_n626), .ZN(new_n967));
  MUX2_X1   g0767(.A(new_n966), .B(new_n663), .S(new_n967), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n751), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n701), .B(KEYINPUT41), .Z(new_n971));
  NAND3_X1  g0771(.A1(new_n523), .A2(new_n686), .A3(new_n682), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n515), .B2(new_n689), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n667), .A2(new_n606), .A3(new_n689), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n682), .B1(new_n584), .B2(new_n588), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n655), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT104), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT104), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n698), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT45), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT44), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n698), .B2(new_n976), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n973), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n694), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n981), .A2(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n694), .A3(new_n984), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n994));
  INV_X1    g0794(.A(new_n693), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n695), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n972), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT105), .A3(new_n688), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n972), .A3(new_n999), .A4(new_n996), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n991), .A2(new_n740), .A3(new_n993), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n971), .B1(new_n1002), .B2(new_n740), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n744), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n696), .A2(new_n976), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n515), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n665), .B1(new_n976), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1008), .B2(new_n689), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n968), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n968), .A2(new_n1011), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n694), .A2(new_n977), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n970), .B1(new_n1004), .B2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n740), .A2(new_n1001), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n998), .B(new_n1000), .C1(new_n731), .C2(new_n739), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n701), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n269), .B1(new_n770), .B2(new_n789), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n767), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1022));
  INV_X1    g0822(.A(G322), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n784), .B2(new_n781), .C1(new_n1023), .C2(new_n788), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n792), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n844), .A2(G294), .B1(G283), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT49), .Z(new_n1031));
  AOI211_X1 g0831(.A(new_n1021), .B(new_n1031), .C1(G116), .C2(new_n840), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n844), .A2(G77), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G68), .A2(new_n832), .B1(new_n771), .B2(G150), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n202), .C2(new_n766), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n269), .B1(new_n840), .B2(G97), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n253), .ZN(new_n1037));
  INV_X1    g0837(.A(G159), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1036), .B1(new_n784), .B2(new_n1037), .C1(new_n1038), .C2(new_n788), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n633), .A2(new_n804), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n759), .B1(new_n1032), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n302), .B1(new_n263), .B2(new_n368), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n703), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT109), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n253), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT50), .B1(new_n253), .B2(new_n202), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n939), .B(new_n1049), .C1(new_n234), .C2(new_n302), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(G107), .B2(new_n212), .C1(new_n703), .C2(new_n753), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n857), .B1(new_n1051), .B2(new_n760), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1042), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n995), .B2(new_n751), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1001), .B2(new_n744), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1020), .A2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n991), .A2(new_n993), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1018), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n701), .A3(new_n1002), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n989), .A2(new_n990), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n694), .B1(new_n992), .B2(new_n984), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT110), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT110), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n991), .A2(new_n993), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n744), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n977), .A2(new_n751), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT111), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n939), .A2(new_n246), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n761), .B1(G97), .B2(new_n700), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n778), .A2(new_n263), .B1(new_n955), .B2(new_n770), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT112), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n788), .A2(new_n835), .B1(new_n1038), .B2(new_n766), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n805), .A2(G77), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n274), .B1(new_n774), .B2(new_n797), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1037), .A2(new_n780), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G50), .C2(new_n783), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G317), .A2(new_n787), .B1(new_n767), .B2(G311), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n780), .A2(new_n790), .B1(new_n770), .B2(new_n1023), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n274), .B(new_n1083), .C1(G107), .C2(new_n840), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G116), .A2(new_n1028), .B1(new_n783), .B2(G303), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n773), .C2(new_n778), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1073), .A2(new_n1080), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n857), .B(new_n1070), .C1(new_n1087), .C2(new_n759), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1067), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1059), .A2(new_n1065), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n743), .B1(new_n1057), .B2(KEYINPUT110), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1093), .A2(new_n1064), .B1(new_n1067), .B2(new_n1088), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(KEYINPUT113), .A3(new_n1059), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(G390));
  NOR2_X1   g0896(.A1(new_n824), .A2(new_n674), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n915), .A2(KEYINPUT114), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1098), .A2(new_n729), .A3(new_n906), .A4(new_n1097), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n737), .A2(new_n682), .A3(new_n822), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n907), .B1(new_n1100), .B2(new_n823), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n872), .B1(new_n356), .B2(new_n865), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n889), .B1(new_n1102), .B2(KEYINPUT38), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1101), .A2(new_n894), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(KEYINPUT101), .B(new_n891), .C1(new_n898), .C2(new_n878), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n900), .B1(new_n899), .B2(KEYINPUT39), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n892), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n827), .A2(new_n823), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n894), .B1(new_n1109), .B2(new_n906), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1099), .B(new_n1105), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n915), .A2(new_n1097), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1112), .A2(KEYINPUT114), .A3(new_n907), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n893), .B2(new_n901), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n1104), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1115), .A3(new_n744), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n858), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n745), .B1(new_n253), .B2(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n269), .B1(new_n263), .B2(new_n774), .C1(new_n788), .C2(new_n773), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G107), .B2(new_n783), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n798), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n766), .A2(new_n535), .B1(new_n780), .B2(new_n538), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G294), .B2(new_n771), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1076), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n953), .A2(new_n783), .B1(new_n787), .B2(G128), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n269), .B1(new_n767), .B2(G132), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n840), .A2(G50), .B1(new_n771), .B2(G125), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT116), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1128), .B1(new_n1038), .B2(new_n804), .C1(new_n780), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n844), .A2(G150), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1118), .B1(new_n1135), .B2(new_n759), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1108), .B2(new_n750), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1116), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n470), .A2(G330), .A3(new_n915), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n654), .A2(new_n911), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n906), .B1(new_n729), .B2(new_n1097), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1112), .A2(new_n907), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1109), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n729), .A2(new_n906), .A3(new_n1097), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1112), .A2(new_n907), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n823), .A3(new_n1100), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT115), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1111), .A2(new_n1115), .A3(new_n1147), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n701), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1138), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  NOR2_X1   g0954(.A1(new_n680), .A2(new_n366), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT55), .Z(new_n1156));
  OR2_X1    g0956(.A1(new_n389), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n389), .A2(new_n1156), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n919), .B1(new_n876), .B2(new_n874), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n915), .A2(new_n916), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT40), .B1(new_n1103), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n674), .B(new_n1164), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(G330), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n910), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1164), .B1(new_n920), .B2(new_n674), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(G330), .A3(new_n1169), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1173), .A2(new_n1174), .B1(new_n902), .B2(new_n909), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n744), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT118), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1164), .A2(new_n749), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n745), .B1(G50), .B2(new_n1117), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n265), .B(new_n301), .C1(new_n774), .C2(new_n807), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  INV_X1    g0981(.A(G137), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n766), .A2(new_n1181), .B1(new_n780), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n784), .A2(new_n842), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G125), .C2(new_n787), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n835), .B2(new_n804), .C1(new_n778), .C2(new_n1131), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1180), .B(new_n1187), .C1(G124), .C2(new_n771), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(KEYINPUT59), .B2(new_n1186), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n784), .A2(new_n538), .B1(new_n788), .B2(new_n535), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n269), .A2(new_n301), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n766), .A2(new_n447), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n774), .A2(new_n250), .B1(new_n770), .B2(new_n773), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n632), .A2(new_n832), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1194), .A2(new_n957), .A3(new_n1033), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1191), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1189), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1179), .B1(new_n1201), .B2(new_n759), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1178), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1176), .A2(new_n1177), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n910), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1173), .A2(new_n902), .A3(new_n1174), .A4(new_n909), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n743), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1203), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT118), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1140), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1151), .A2(new_n1211), .B1(new_n1206), .B2(new_n1205), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n701), .B1(new_n1212), .B2(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1151), .A2(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1214), .A2(KEYINPUT57), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1213), .B2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n907), .A2(new_n749), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n745), .B1(G68), .B2(new_n1117), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n780), .A2(new_n835), .B1(new_n770), .B2(new_n1181), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n274), .B1(new_n250), .B2(new_n774), .C1(new_n788), .C2(new_n842), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n767), .C2(new_n953), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n844), .A2(G159), .B1(new_n1130), .B2(new_n783), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n202), .C2(new_n804), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n778), .A2(new_n538), .B1(new_n527), .B2(new_n770), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT120), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n767), .A2(G283), .B1(new_n832), .B2(G107), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n784), .B2(new_n535), .C1(new_n790), .C2(new_n788), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n269), .B1(new_n774), .B2(new_n368), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT119), .ZN(new_n1231));
  OR3_X1    g1031(.A1(new_n1229), .A2(new_n1040), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1225), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1220), .B1(new_n1233), .B2(new_n759), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1218), .A2(new_n744), .B1(new_n1219), .B2(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1147), .A2(new_n971), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1218), .A2(new_n1211), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  NAND3_X1  g1038(.A1(new_n1020), .A2(new_n817), .A3(new_n1055), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1239), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G390), .A2(new_n1240), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1041(.A(G375), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n678), .A2(G343), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT121), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT122), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1153), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G407), .A2(G213), .A3(new_n1246), .ZN(G409));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT113), .B1(new_n1094), .B2(new_n1059), .ZN(new_n1249));
  AND4_X1   g1049(.A1(KEYINPUT113), .A2(new_n1059), .A3(new_n1065), .A4(new_n1089), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT123), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G387), .A2(new_n1239), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1092), .A2(new_n1095), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1239), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n970), .C1(new_n1004), .C2(new_n1016), .ZN(new_n1257));
  AND4_X1   g1057(.A1(new_n1251), .A2(new_n1253), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1251), .A2(new_n1255), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1248), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n971), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1152), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1138), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(G375), .B2(new_n1153), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1244), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1147), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1237), .B1(KEYINPUT60), .B2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1143), .A2(new_n1146), .A3(KEYINPUT60), .A4(new_n1140), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n701), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1235), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n860), .A3(new_n831), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G384), .B(new_n1235), .C1(new_n1272), .C2(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G2897), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1244), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1245), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1260), .B1(new_n1270), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1269), .A2(new_n1244), .A3(new_n1279), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1269), .A2(new_n1283), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1278), .A2(new_n1288), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1286), .B(new_n1289), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1248), .B1(new_n1296), .B2(new_n1290), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1278), .A2(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1269), .A2(new_n1283), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(new_n1298), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1287), .A2(KEYINPUT125), .A3(new_n1298), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1297), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1295), .B1(new_n1305), .B2(new_n1307), .ZN(G405));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(G375), .B2(new_n1153), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(G378), .B2(new_n1242), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G375), .A2(new_n1309), .A3(new_n1153), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1307), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1306), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(G402));
endmodule


