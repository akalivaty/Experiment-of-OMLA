//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT77), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n210), .A2(new_n219), .A3(new_n216), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR3_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n207), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT78), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(KEYINPUT78), .C2(new_n214), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n225), .A2(new_n228), .A3(new_n209), .A4(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n221), .A2(KEYINPUT80), .A3(new_n229), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT16), .A3(new_n235), .ZN(new_n236));
  OAI221_X1 g035(.A(new_n236), .B1(KEYINPUT81), .B2(G8gat), .C1(new_n235), .C2(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n232), .A2(new_n241), .A3(new_n233), .ZN(new_n242));
  INV_X1    g041(.A(new_n239), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n229), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n202), .B(new_n240), .C1(new_n242), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n243), .B(new_n244), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n240), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n202), .B(KEYINPUT13), .Z(new_n252));
  INV_X1    g051(.A(new_n240), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n239), .B1(new_n232), .B2(new_n233), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n248), .A2(new_n261), .A3(new_n251), .A4(new_n255), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n267));
  XOR2_X1   g066(.A(G141gat), .B(G148gat), .Z(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(KEYINPUT2), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G141gat), .B(G148gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n272), .B(new_n271), .C1(new_n276), .C2(KEYINPUT2), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT70), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n275), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT1), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n284), .B(new_n286), .C1(new_n282), .C2(KEYINPUT1), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n275), .A2(new_n277), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(KEYINPUT3), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n290), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT4), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n293), .A2(new_n294), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n279), .A2(new_n280), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  INV_X1    g102(.A(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n267), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n300), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n278), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n291), .B1(new_n311), .B2(KEYINPUT3), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT5), .B1(new_n313), .B2(new_n294), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT71), .B(KEYINPUT0), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n307), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n306), .B2(new_n314), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  AND2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(KEYINPUT22), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT67), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  INV_X1    g144(.A(G169gat), .ZN(new_n346));
  INV_X1    g145(.A(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n348), .A2(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n344), .A2(new_n350), .A3(KEYINPUT25), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OR3_X1    g154(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(new_n346), .C2(new_n347), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n359), .A2(KEYINPUT28), .A3(new_n342), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT28), .B1(new_n359), .B2(new_n342), .ZN(new_n361));
  OAI221_X1 g160(.A(new_n358), .B1(new_n341), .B2(new_n342), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n337), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n368), .A3(new_n337), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n334), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n336), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n364), .A2(new_n368), .A3(new_n366), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n337), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n371), .B(new_n374), .C1(new_n378), .C2(new_n334), .ZN(new_n379));
  NOR4_X1   g178(.A1(new_n306), .A2(new_n314), .A3(new_n323), .A4(new_n320), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n325), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n355), .A2(new_n362), .A3(new_n365), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n365), .B1(new_n355), .B2(new_n362), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n336), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n333), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT29), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n375), .B1(new_n388), .B2(new_n336), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n333), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n374), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n333), .B1(new_n367), .B2(new_n370), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(KEYINPUT37), .C1(new_n378), .C2(new_n333), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT38), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n371), .B1(new_n378), .B2(new_n334), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(KEYINPUT37), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n395), .A2(new_n396), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n311), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n368), .B1(new_n290), .B2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n333), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n401), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n290), .B2(new_n403), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  OR3_X1    g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT73), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n410), .B1(new_n407), .B2(new_n409), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n411), .A2(new_n418), .B1(new_n416), .B2(new_n415), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT69), .B1(new_n379), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n390), .A2(new_n425), .A3(KEYINPUT30), .A4(new_n374), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n379), .A2(new_n423), .ZN(new_n427));
  INV_X1    g226(.A(new_n374), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n397), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n424), .A2(new_n426), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n313), .A2(new_n433), .A3(new_n294), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT75), .B1(new_n435), .B2(new_n304), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n313), .B2(new_n294), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n304), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n303), .A2(new_n304), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n438), .A2(KEYINPUT39), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n441), .A3(new_n320), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT40), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT40), .A4(new_n320), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n322), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n422), .B1(new_n431), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n400), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n424), .A2(new_n427), .A3(new_n429), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n306), .A2(new_n314), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n321), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n325), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n449), .A2(new_n450), .A3(new_n453), .A4(new_n426), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT6), .B1(new_n451), .B2(new_n321), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n380), .B1(new_n455), .B2(new_n324), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT72), .B1(new_n430), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n422), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n363), .A2(new_n296), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n355), .A2(new_n362), .A3(new_n288), .A4(new_n289), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n459), .A2(G227gat), .A3(G233gat), .A4(new_n460), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G15gat), .B(G43gat), .Z(new_n472));
  XNOR2_X1  g271(.A(G71gat), .B(G99gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n474), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n468), .B(KEYINPUT32), .C1(new_n470), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n467), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n467), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n479), .A2(new_n480), .B1(new_n464), .B2(new_n463), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n477), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n466), .A3(new_n465), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n464), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n478), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n481), .A2(new_n485), .A3(new_n487), .A4(KEYINPUT36), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n448), .A2(new_n458), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n421), .B1(new_n481), .B2(new_n485), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n454), .A2(new_n457), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n325), .B1(new_n381), .B2(new_n382), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(new_n431), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n266), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT9), .ZN(new_n503));
  NAND2_X1  g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  INV_X1    g305(.A(G57gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT83), .A2(G57gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(G64gat), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G64gat), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT84), .B1(new_n511), .B2(G57gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(KEYINPUT84), .A3(G64gat), .A4(new_n509), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n513), .A2(KEYINPUT85), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT85), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n502), .B1(KEYINPUT82), .B2(new_n504), .ZN(new_n518));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(KEYINPUT82), .A2(KEYINPUT9), .ZN(new_n520));
  OAI221_X1 g319(.A(new_n518), .B1(KEYINPUT82), .B2(new_n504), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G127gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n243), .B1(new_n523), .B2(new_n522), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT86), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G155gat), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT88), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n531), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n531), .B2(new_n532), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G99gat), .ZN(new_n548));
  INV_X1    g347(.A(G106gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT8), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n249), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n244), .B(new_n561), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n569));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n572), .A3(new_n565), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n568), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n543), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n517), .A2(new_n521), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n557), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n557), .A2(new_n517), .A3(new_n521), .A4(new_n579), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n522), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n558), .A3(KEYINPUT10), .A4(new_n560), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT93), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n582), .B2(new_n584), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n592), .A2(new_n600), .A3(new_n594), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n597), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n590), .B1(new_n585), .B2(new_n587), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT95), .B(new_n603), .C1(new_n604), .C2(new_n593), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT96), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(KEYINPUT96), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n578), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n501), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n453), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT97), .B(G1gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(G1324gat));
  NAND3_X1  g417(.A1(new_n501), .A2(new_n430), .A3(new_n614), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT16), .B(G8gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n621), .A2(KEYINPUT42), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(KEYINPUT42), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(G8gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(G1325gat));
  INV_X1    g424(.A(new_n492), .ZN(new_n626));
  OAI21_X1  g425(.A(G15gat), .B1(new_n615), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n486), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(G15gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n615), .B2(new_n629), .ZN(G1326gat));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n422), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT98), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT43), .B(G22gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1327gat));
  AND3_X1   g433(.A1(new_n602), .A2(KEYINPUT96), .A3(new_n609), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n610), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n542), .A2(new_n636), .A3(new_n576), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT99), .Z(new_n638));
  NAND4_X1  g437(.A1(new_n501), .A2(new_n638), .A3(new_n204), .A4(new_n456), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT45), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n448), .A2(new_n458), .A3(new_n492), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n500), .A2(KEYINPUT101), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n496), .A2(new_n643), .A3(new_n499), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n577), .A2(KEYINPUT44), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT102), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n644), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n643), .B1(new_n496), .B2(new_n499), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n493), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n646), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n493), .A2(new_n500), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n576), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n648), .A2(new_n653), .B1(KEYINPUT44), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n613), .B(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n265), .A3(new_n542), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n656), .A2(new_n453), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n640), .B1(new_n659), .B2(new_n204), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n648), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(KEYINPUT44), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n205), .B1(new_n664), .B2(new_n430), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n501), .A2(new_n205), .A3(new_n430), .A4(new_n638), .ZN(new_n666));
  NAND2_X1  g465(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n661), .B1(new_n665), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n656), .A2(new_n431), .A3(new_n658), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n674), .B(KEYINPUT104), .C1(new_n675), .C2(new_n205), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(G1329gat));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n663), .ZN(new_n678));
  INV_X1    g477(.A(new_n658), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n626), .A2(new_n213), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n501), .A2(new_n486), .A3(new_n638), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n682), .A2(new_n213), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT106), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n681), .B2(new_n683), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(G1330gat));
  NOR2_X1   g487(.A1(new_n422), .A2(G50gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n501), .A2(new_n638), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT108), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n678), .A2(new_n421), .A3(new_n679), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(G50gat), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n694));
  AOI21_X1  g493(.A(new_n211), .B1(new_n664), .B2(new_n421), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(KEYINPUT48), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n693), .A2(new_n694), .B1(new_n695), .B2(new_n696), .ZN(G1331gat));
  NOR4_X1   g496(.A1(new_n645), .A2(new_n265), .A3(new_n578), .A4(new_n657), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n456), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n508), .A2(new_n509), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1332gat));
  XNOR2_X1  g500(.A(new_n430), .B(KEYINPUT109), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT49), .B(G64gat), .Z(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(G1333gat));
  NAND2_X1  g506(.A1(new_n698), .A2(new_n492), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n628), .A2(G71gat), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(G71gat), .B1(new_n698), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g510(.A1(new_n698), .A2(new_n421), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G78gat), .ZN(G1335gat));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT51), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n543), .A2(new_n265), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n577), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n645), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n645), .B2(new_n719), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n613), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n545), .A3(new_n456), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n717), .A2(new_n613), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n662), .B2(new_n663), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727), .B2(new_n453), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1336gat));
  INV_X1    g528(.A(new_n657), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n702), .A2(G92gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n720), .A2(new_n730), .A3(new_n721), .A4(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n725), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n678), .A2(new_n430), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n544), .A2(new_n546), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n726), .A2(new_n703), .B1(new_n544), .B2(new_n546), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n741), .ZN(G1337gat));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n548), .A3(new_n486), .ZN(new_n743));
  OAI21_X1  g542(.A(G99gat), .B1(new_n727), .B2(new_n626), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1338gat));
  AOI21_X1  g544(.A(new_n549), .B1(new_n726), .B2(new_n421), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n422), .A2(G106gat), .ZN(new_n747));
  AND4_X1   g546(.A1(new_n730), .A2(new_n720), .A3(new_n721), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT53), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n656), .A2(new_n422), .A3(new_n725), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n750), .B(new_n751), .C1(new_n752), .C2(new_n549), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(G1339gat));
  AOI21_X1  g553(.A(new_n202), .B1(new_n250), .B2(new_n240), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n253), .A2(new_n254), .A3(new_n252), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n260), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n264), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n635), .B2(new_n610), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n585), .A2(new_n590), .A3(new_n587), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n592), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n597), .B1(new_n604), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n763), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n265), .A2(new_n602), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n576), .B1(new_n759), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n602), .A2(new_n764), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n576), .A2(new_n758), .A3(new_n770), .A4(new_n767), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n542), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n543), .A2(new_n266), .A3(new_n577), .A4(new_n636), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n494), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n703), .A2(new_n453), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n265), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G113gat), .ZN(G1340gat));
  AND3_X1   g581(.A1(new_n780), .A2(G120gat), .A3(new_n730), .ZN(new_n783));
  AOI21_X1  g582(.A(G120gat), .B1(new_n780), .B2(new_n613), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1341gat));
  NAND2_X1  g584(.A1(new_n780), .A2(new_n543), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g586(.A1(new_n576), .A2(new_n456), .A3(new_n431), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(G134gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT56), .Z(new_n791));
  OAI21_X1  g590(.A(G134gat), .B1(new_n779), .B2(new_n577), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1343gat));
  AOI21_X1  g592(.A(new_n422), .B1(new_n772), .B2(new_n773), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n626), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n266), .A2(G141gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(KEYINPUT114), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n795), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g602(.A1(new_n265), .A2(new_n602), .A3(new_n764), .A4(new_n767), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n759), .B2(KEYINPUT112), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n613), .A2(new_n806), .A3(new_n758), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n576), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n542), .B1(new_n808), .B2(new_n771), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n422), .B1(new_n809), .B2(new_n773), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n265), .B(new_n803), .C1(new_n810), .C2(new_n802), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G141gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n800), .A2(KEYINPUT114), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n801), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n800), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(KEYINPUT58), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n799), .B1(new_n811), .B2(G141gat), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(KEYINPUT113), .A3(new_n813), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n815), .B1(new_n818), .B2(new_n820), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n794), .A2(KEYINPUT57), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n810), .B2(KEYINPUT57), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n613), .A3(new_n796), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n825));
  INV_X1    g624(.A(G148gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n613), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n803), .ZN(new_n828));
  INV_X1    g627(.A(new_n810), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(KEYINPUT57), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n830), .B2(new_n613), .ZN(new_n831));
  OAI221_X1 g630(.A(new_n825), .B1(new_n797), .B2(new_n827), .C1(new_n831), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g631(.A(new_n269), .B1(new_n830), .B2(new_n543), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n797), .A2(G155gat), .A3(new_n542), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(new_n834), .ZN(G1346gat));
  OAI211_X1 g634(.A(new_n576), .B(new_n803), .C1(new_n810), .C2(new_n802), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n270), .B1(new_n836), .B2(KEYINPUT115), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(KEYINPUT115), .B2(new_n836), .ZN(new_n838));
  INV_X1    g637(.A(new_n794), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n492), .A2(G162gat), .A3(new_n788), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G1347gat));
  NOR3_X1   g640(.A1(new_n628), .A2(new_n456), .A3(new_n431), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n422), .B1(new_n842), .B2(KEYINPUT118), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(KEYINPUT118), .B2(new_n842), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n774), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n346), .A3(new_n266), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n703), .B2(new_n494), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n702), .A2(new_n776), .A3(KEYINPUT116), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n453), .A3(new_n774), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n265), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n846), .B1(new_n854), .B2(new_n346), .ZN(G1348gat));
  NOR3_X1   g654(.A1(new_n845), .A2(new_n347), .A3(new_n657), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n613), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n347), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n347), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(G1349gat));
  INV_X1    g661(.A(new_n845), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n341), .B1(new_n863), .B2(new_n543), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(KEYINPUT60), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n775), .A2(new_n456), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(new_n359), .A3(new_n543), .A4(new_n850), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n865), .A2(KEYINPUT60), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(G1350gat));
  NAND4_X1  g670(.A1(new_n852), .A2(new_n342), .A3(new_n576), .A4(new_n853), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G190gat), .B1(new_n845), .B2(new_n577), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT61), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1351gat));
  INV_X1    g676(.A(G197gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n431), .A2(new_n456), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n626), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT124), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n823), .A2(new_n265), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(KEYINPUT125), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(KEYINPUT125), .B2(new_n882), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n626), .A2(new_n421), .A3(new_n703), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n867), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G197gat), .A3(new_n266), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n890), .ZN(G1352gat));
  OR3_X1    g690(.A1(new_n887), .A2(G204gat), .A3(new_n636), .ZN(new_n892));
  AND2_X1   g691(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n893));
  NOR2_X1   g692(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n823), .A2(new_n730), .A3(new_n881), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G204gat), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n895), .B(new_n897), .C1(new_n893), .C2(new_n892), .ZN(G1353gat));
  NOR3_X1   g697(.A1(new_n887), .A2(G211gat), .A3(new_n542), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT127), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n901));
  INV_X1    g700(.A(new_n823), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n626), .A2(new_n543), .A3(new_n879), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(G211gat), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G211gat), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT63), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n900), .A2(new_n904), .A3(new_n906), .ZN(G1354gat));
  AND3_X1   g706(.A1(new_n823), .A2(new_n576), .A3(new_n881), .ZN(new_n908));
  INV_X1    g707(.A(G218gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n576), .A2(new_n909), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n908), .A2(new_n909), .B1(new_n887), .B2(new_n910), .ZN(G1355gat));
endmodule


