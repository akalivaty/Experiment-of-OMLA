//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(G116), .B(G119), .Z(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT2), .B(G113), .Z(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT66), .B1(new_n195), .B2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT66), .B(new_n198), .C1(new_n195), .C2(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G131), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n203), .A3(new_n199), .A4(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT0), .B(G128), .Z(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT65), .A2(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(G143), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n206), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(G143), .A3(new_n210), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(KEYINPUT0), .A3(G128), .A4(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(new_n215), .A3(G128), .A4(new_n217), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n210), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT65), .A2(G146), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n224), .A2(new_n225), .A3(new_n216), .ZN(new_n226));
  OAI21_X1  g040(.A(G128), .B1(new_n226), .B2(new_n221), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n224), .A2(new_n225), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n212), .B1(new_n229), .B2(G143), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n215), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT65), .B(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n213), .B1(new_n235), .B2(new_n216), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT70), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n223), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n239), .B2(G134), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n195), .A3(G137), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(new_n242), .C1(new_n195), .C2(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT68), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n246), .A3(G131), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n204), .A3(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT30), .B(new_n220), .C1(new_n238), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n214), .A2(new_n218), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n202), .B2(new_n204), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n228), .B1(new_n227), .B2(new_n230), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT70), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n222), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n245), .A2(new_n204), .A3(new_n247), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n194), .B(new_n249), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G210), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n261), .B(KEYINPUT27), .Z(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  XNOR2_X1  g078(.A(new_n194), .B(KEYINPUT71), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(new_n220), .C1(new_n238), .C2(new_n248), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT31), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n220), .A4(new_n265), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n194), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n270), .B2(new_n220), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n264), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n269), .B2(new_n272), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n280), .A2(new_n281), .A3(new_n264), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n268), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n258), .A2(new_n284), .A3(new_n264), .A4(new_n266), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT72), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n278), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n281), .B1(new_n280), .B2(new_n264), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n289), .A2(new_n290), .B1(KEYINPUT31), .B2(new_n267), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n285), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n187), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n256), .A2(new_n265), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n273), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n258), .A2(new_n266), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n278), .ZN(new_n307));
  AOI211_X1 g121(.A(KEYINPUT76), .B(new_n264), .C1(new_n258), .C2(new_n266), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n280), .B2(new_n264), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n299), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n278), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n306), .A2(new_n305), .A3(new_n278), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n310), .ZN(new_n317));
  INV_X1    g131(.A(new_n304), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT77), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT32), .B(new_n187), .C1(new_n283), .C2(new_n286), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n298), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G234), .ZN(new_n324));
  OAI21_X1  g138(.A(G217), .B1(new_n324), .B2(G902), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT78), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT79), .B1(new_n232), .B2(G119), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G119), .B(G128), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  AOI22_X1  g145(.A1(new_n329), .A2(G110), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n335), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G146), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n208), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n329), .A2(G110), .B1(new_n330), .B2(new_n331), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(G146), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n229), .A2(new_n333), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(new_n345), .A3(KEYINPUT81), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n345), .A3(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n348), .B(KEYINPUT80), .Z(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n341), .B2(new_n345), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n349), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n355), .A2(new_n300), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n355), .B2(new_n300), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n326), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n326), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  OAI21_X1  g179(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n369), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n370), .A2(new_n373), .A3(new_n377), .A4(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n381), .A3(G101), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n214), .A2(new_n382), .A3(new_n218), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n368), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n219), .A2(new_n379), .A3(KEYINPUT83), .A4(new_n382), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n369), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n372), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n232), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n215), .B2(new_n217), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n223), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n384), .A2(new_n385), .B1(new_n386), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n254), .A2(KEYINPUT10), .A3(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n205), .ZN(new_n398));
  INV_X1    g212(.A(new_n205), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n260), .A2(G227), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT85), .A2(KEYINPUT12), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n238), .A2(new_n410), .A3(new_n390), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n205), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n223), .B(new_n391), .C1(new_n231), .C2(new_n237), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n394), .A2(KEYINPUT84), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n406), .B(new_n409), .C1(new_n412), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n399), .B1(new_n413), .B2(new_n410), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT84), .B(new_n394), .C1(new_n254), .C2(new_n391), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n407), .A4(new_n408), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(KEYINPUT87), .ZN(new_n420));
  INV_X1    g234(.A(new_n404), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n400), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT87), .B1(new_n416), .B2(new_n419), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n405), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT86), .B(G469), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n300), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n398), .A2(new_n400), .A3(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n416), .A2(new_n419), .A3(new_n400), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n404), .ZN(new_n430));
  OAI21_X1  g244(.A(G469), .B1(new_n430), .B2(G902), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n367), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(G234), .A2(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(G952), .A3(new_n260), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(G902), .A3(G953), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n379), .A2(new_n194), .A3(new_n382), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n192), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g258(.A(G116), .ZN(new_n445));
  OR3_X1    g259(.A1(new_n445), .A2(KEYINPUT5), .A3(G119), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(G113), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n391), .A2(new_n193), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT6), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n448), .ZN(new_n451));
  INV_X1    g265(.A(new_n443), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n450), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n219), .A2(G125), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n238), .B2(G125), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI221_X1 g273(.A(new_n455), .B1(new_n457), .B2(G953), .C1(new_n238), .C2(G125), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n459), .B(new_n460), .C1(KEYINPUT7), .C2(new_n458), .ZN(new_n464));
  OR3_X1    g278(.A1(new_n456), .A2(KEYINPUT7), .A3(new_n458), .ZN(new_n465));
  INV_X1    g279(.A(new_n449), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n193), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n390), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n448), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n443), .B(KEYINPUT8), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n462), .A2(new_n463), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n463), .B1(new_n462), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n433), .B(new_n441), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n476));
  NOR2_X1   g290(.A1(KEYINPUT88), .A2(G143), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  OR2_X1    g293(.A1(KEYINPUT88), .A2(G143), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n476), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n203), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT89), .B1(new_n483), .B2(KEYINPUT17), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n339), .A2(new_n340), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n479), .A2(new_n482), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(KEYINPUT17), .A3(G131), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n484), .A2(new_n485), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n369), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n481), .B1(new_n493), .B2(new_n203), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n478), .A2(KEYINPUT18), .A3(G131), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n344), .B1(new_n208), .B2(new_n333), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n490), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n492), .B1(new_n490), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n300), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT90), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(new_n300), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(G475), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n490), .A2(new_n492), .A3(new_n497), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n333), .B(KEYINPUT19), .Z(new_n506));
  OAI211_X1 g320(.A(new_n483), .B(new_n343), .C1(new_n235), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  INV_X1    g322(.A(new_n492), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G475), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n300), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n511), .A2(new_n516), .A3(new_n513), .A4(new_n300), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT13), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n232), .A2(KEYINPUT13), .A3(G143), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n195), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n520), .A2(new_n522), .B1(new_n195), .B2(new_n519), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT91), .B(G122), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n445), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n445), .B2(G122), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n372), .ZN(new_n527));
  AOI211_X1 g341(.A(G107), .B(new_n525), .C1(new_n445), .C2(G122), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n372), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n445), .A2(G122), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g346(.A(G107), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n519), .B(new_n195), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n365), .A2(new_n537), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n529), .A2(new_n535), .A3(new_n538), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n542), .A2(KEYINPUT15), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n545));
  AOI211_X1 g359(.A(G902), .B(new_n545), .C1(new_n540), .C2(new_n541), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n504), .A2(new_n518), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n475), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n432), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n323), .A2(new_n364), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(G101), .ZN(G3));
  AND2_X1   g366(.A1(new_n288), .A2(new_n296), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n291), .B2(new_n293), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n312), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n300), .B1(new_n283), .B2(new_n286), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT92), .A3(G472), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n367), .B(new_n363), .C1(new_n427), .C2(new_n431), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n504), .A2(new_n518), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n540), .A2(new_n541), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT33), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n540), .A2(new_n565), .A3(new_n541), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(G478), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n543), .A2(new_n300), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n542), .B2(new_n543), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n440), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n462), .A2(new_n472), .ZN(new_n574));
  INV_X1    g388(.A(new_n463), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n462), .A2(new_n463), .A3(new_n472), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT93), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n433), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n561), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT34), .B(G104), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G6));
  INV_X1    g398(.A(new_n547), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n504), .A3(new_n518), .A4(new_n441), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT94), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n561), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G107), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G9));
  INV_X1    g404(.A(new_n353), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n341), .A2(new_n345), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n361), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n360), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n550), .A2(new_n553), .A3(new_n559), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT37), .B(G110), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G12));
  NAND2_X1  g413(.A1(new_n432), .A2(new_n596), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n437), .A2(G900), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n435), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n562), .A2(new_n547), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n323), .A2(new_n606), .A3(new_n581), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G128), .ZN(G30));
  INV_X1    g422(.A(new_n267), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n264), .B1(new_n301), .B2(new_n266), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n300), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n298), .A2(new_n322), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n602), .B(KEYINPUT39), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n432), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n576), .A2(new_n577), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n433), .B1(new_n544), .B2(new_n546), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n504), .B2(new_n518), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n623), .A2(new_n360), .A3(new_n595), .A4(new_n625), .ZN(new_n626));
  NOR4_X1   g440(.A1(new_n614), .A2(new_n618), .A3(new_n619), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n216), .ZN(G45));
  AOI211_X1 g443(.A(new_n603), .B(new_n570), .C1(new_n504), .C2(new_n518), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n432), .A2(new_n596), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n323), .A2(new_n581), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n323), .A2(new_n631), .A3(KEYINPUT99), .A4(new_n581), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G146), .ZN(G48));
  AND2_X1   g451(.A1(new_n425), .A2(new_n300), .ZN(new_n638));
  INV_X1    g452(.A(G469), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n366), .B(new_n427), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n580), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n323), .A2(new_n364), .A3(new_n573), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT41), .B(G113), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G15));
  NAND4_X1  g459(.A1(new_n323), .A2(new_n364), .A3(new_n587), .A4(new_n641), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G116), .ZN(G18));
  AND2_X1   g461(.A1(new_n504), .A2(new_n518), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(new_n596), .A3(new_n547), .A4(new_n441), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n640), .A2(new_n580), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n323), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G119), .ZN(G21));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(G472), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n557), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n302), .A2(new_n278), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n268), .A3(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n293), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT101), .B1(new_n655), .B2(new_n268), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n187), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n360), .A2(KEYINPUT103), .A3(new_n362), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT103), .B1(new_n360), .B2(new_n362), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n625), .B(new_n441), .C1(new_n578), .C2(new_n579), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  AND3_X1   g482(.A1(new_n654), .A2(new_n596), .A3(new_n659), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n641), .A2(new_n669), .A3(new_n630), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G125), .ZN(G27));
  INV_X1    g485(.A(new_n663), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT32), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n287), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n319), .A2(KEYINPUT77), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n299), .B(new_n312), .C1(new_n317), .C2(new_n318), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n322), .A2(KEYINPUT105), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n294), .A2(new_n679), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n672), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n576), .A2(new_n577), .A3(new_n433), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n429), .A2(new_n404), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n398), .A2(new_n400), .A3(new_n421), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n398), .A2(KEYINPUT104), .A3(new_n400), .A4(new_n421), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n300), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n367), .B(new_n683), .C1(new_n691), .C2(new_n427), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n630), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT42), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n572), .A2(KEYINPUT42), .A3(new_n603), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n323), .A2(new_n364), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n694), .A2(KEYINPUT106), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT106), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G131), .ZN(G33));
  NAND2_X1  g514(.A1(new_n323), .A2(new_n364), .ZN(new_n701));
  INV_X1    g515(.A(new_n683), .ZN(new_n702));
  INV_X1    g516(.A(new_n427), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n639), .B1(new_n689), .B2(new_n300), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n366), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n701), .A2(new_n605), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n195), .ZN(G36));
  NAND2_X1  g521(.A1(new_n648), .A2(new_n571), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT43), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n553), .A2(new_n559), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n596), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n430), .B2(KEYINPUT45), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n689), .A2(new_n715), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n714), .A2(new_n716), .B1(new_n639), .B2(new_n300), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n703), .B1(new_n717), .B2(new_n718), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n367), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n721), .A2(new_n615), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n683), .B1(new_n711), .B2(new_n712), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n713), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n239), .ZN(G39));
  XOR2_X1   g539(.A(new_n721), .B(KEYINPUT47), .Z(new_n726));
  NAND3_X1  g540(.A1(new_n630), .A2(new_n363), .A3(new_n702), .ZN(new_n727));
  OR3_X1    g541(.A1(new_n726), .A2(new_n323), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G140), .ZN(G42));
  NOR2_X1   g543(.A1(new_n638), .A2(new_n639), .ZN(new_n730));
  OR3_X1    g544(.A1(new_n730), .A2(KEYINPUT49), .A3(new_n703), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT49), .B1(new_n730), .B2(new_n703), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n672), .A2(new_n366), .A3(new_n433), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n623), .A3(new_n708), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n614), .A2(new_n731), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n607), .A2(new_n670), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n634), .B2(new_n635), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n625), .B1(new_n578), .B2(new_n579), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n367), .B1(new_n691), .B2(new_n427), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n596), .A2(new_n603), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n613), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n737), .ZN(new_n745));
  AND4_X1   g559(.A1(KEYINPUT52), .A2(new_n636), .A3(new_n745), .A4(new_n743), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n697), .A2(new_n698), .A3(new_n706), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n669), .A2(new_n692), .A3(KEYINPUT108), .A4(new_n630), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n654), .A2(new_n630), .A3(new_n659), .A4(new_n596), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(new_n705), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n702), .A2(new_n648), .A3(new_n547), .A4(new_n602), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n600), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n749), .A2(new_n752), .B1(new_n323), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n648), .A2(new_n585), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n475), .B1(new_n756), .B2(new_n572), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n553), .A2(new_n559), .A3(new_n757), .A4(new_n560), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n597), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n759), .A3(new_n551), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n323), .A2(new_n650), .B1(new_n664), .B2(new_n666), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n642), .A3(new_n646), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n642), .A3(new_n646), .A4(KEYINPUT107), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n748), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n736), .B1(new_n747), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n636), .A2(new_n745), .A3(new_n743), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n738), .A2(KEYINPUT52), .A3(new_n743), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT109), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n744), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n706), .A2(new_n736), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n694), .A2(new_n696), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n776), .A2(new_n760), .A3(new_n777), .A4(new_n762), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n780));
  NAND3_X1  g594(.A1(new_n768), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n775), .A3(new_n773), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT53), .B1(new_n747), .B2(new_n767), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n640), .A2(new_n363), .A3(new_n435), .A4(new_n683), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n614), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n562), .A3(new_n571), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n709), .A2(new_n436), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n640), .A3(new_n683), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n669), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n709), .A2(new_n436), .A3(new_n664), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n795), .A2(new_n433), .A3(new_n623), .A4(new_n640), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n367), .B(new_n427), .C1(new_n638), .C2(new_n639), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n683), .B(new_n795), .C1(new_n726), .C2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n788), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n260), .A2(G952), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n795), .A2(new_n580), .A3(new_n640), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n802), .B1(new_n803), .B2(KEYINPUT113), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(KEYINPUT113), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n790), .A2(new_n572), .ZN(new_n806));
  INV_X1    g620(.A(new_n682), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n793), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT48), .Z(new_n809));
  NOR3_X1   g623(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n801), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n797), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT112), .Z(new_n815));
  NOR2_X1   g629(.A1(new_n800), .A2(new_n788), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n787), .B(new_n811), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(G952), .A2(G953), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n735), .B1(new_n817), .B2(new_n818), .ZN(G75));
  NOR2_X1   g633(.A1(new_n260), .A2(G952), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT116), .Z(new_n821));
  AOI21_X1  g635(.A(new_n300), .B1(new_n768), .B2(new_n779), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n822), .B2(G210), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n823), .B2(KEYINPUT115), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n454), .B(KEYINPUT114), .Z(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT55), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n461), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n828), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n824), .B1(new_n829), .B2(new_n830), .ZN(G51));
  NAND2_X1  g645(.A1(new_n768), .A2(new_n779), .ZN(new_n832));
  INV_X1    g646(.A(new_n780), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n781), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n639), .A2(new_n300), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT57), .Z(new_n838));
  OAI21_X1  g652(.A(new_n425), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n714), .A2(new_n716), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n822), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n820), .B1(new_n839), .B2(new_n841), .ZN(G54));
  NAND3_X1  g656(.A1(new_n822), .A2(KEYINPUT58), .A3(G475), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n820), .B1(new_n843), .B2(new_n512), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n512), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(KEYINPUT117), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(KEYINPUT117), .B2(new_n845), .ZN(G60));
  AND2_X1   g661(.A1(new_n564), .A2(new_n566), .ZN(new_n848));
  INV_X1    g662(.A(new_n787), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n568), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n821), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(new_n852), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n768), .A2(new_n779), .A3(new_n780), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n780), .B1(new_n768), .B2(new_n779), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n862), .B2(KEYINPUT120), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n864), .B(new_n854), .C1(new_n860), .C2(new_n861), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT121), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT119), .B1(new_n835), .B2(new_n855), .ZN(new_n867));
  INV_X1    g681(.A(new_n861), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n821), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n864), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n862), .A2(KEYINPUT120), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n853), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(G63));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT60), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n594), .B(KEYINPUT122), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n832), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT123), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n355), .B1(new_n832), .B2(new_n876), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n854), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g696(.A(G953), .B1(new_n439), .B2(new_n457), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n759), .A2(new_n551), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n764), .B2(new_n765), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n826), .B1(G898), .B2(new_n260), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(G69));
  AOI21_X1  g702(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n724), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n738), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT124), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n722), .A2(new_n807), .A3(new_n740), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n893), .A2(new_n728), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n748), .B(KEYINPUT125), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n260), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(new_n506), .Z(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(G900), .B2(G953), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n683), .B1(new_n756), .B2(new_n572), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n432), .A3(new_n615), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n728), .B(new_n891), .C1(new_n701), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n905));
  INV_X1    g719(.A(new_n738), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n628), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n628), .B2(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n899), .B1(new_n909), .B2(G953), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n901), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n901), .B2(new_n910), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n890), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n901), .A2(new_n910), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n889), .A3(new_n912), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G72));
  XNOR2_X1  g733(.A(new_n306), .B(KEYINPUT127), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n895), .A2(new_n885), .A3(new_n896), .ZN(new_n921));
  NAND2_X1  g735(.A1(G472), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT63), .Z(new_n923));
  AOI211_X1 g737(.A(new_n264), .B(new_n920), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n923), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n909), .B2(new_n885), .ZN(new_n926));
  INV_X1    g740(.A(new_n920), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n278), .A3(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n925), .B(new_n785), .C1(new_n309), .C2(new_n267), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n924), .A2(new_n928), .A3(new_n820), .A4(new_n929), .ZN(G57));
endmodule


