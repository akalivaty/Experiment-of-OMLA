

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  NOR2_X1 U324 ( .A1(n527), .A2(n460), .ZN(n485) );
  XNOR2_X1 U325 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U326 ( .A(n465), .B(KEYINPUT99), .ZN(n556) );
  XNOR2_X1 U327 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n429) );
  XNOR2_X1 U328 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U329 ( .A(KEYINPUT36), .B(n549), .Z(n476) );
  XNOR2_X1 U330 ( .A(n461), .B(KEYINPUT125), .ZN(n586) );
  XNOR2_X1 U331 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U332 ( .A(n309), .B(n308), .Z(n292) );
  XOR2_X1 U333 ( .A(n410), .B(KEYINPUT73), .Z(n293) );
  AND2_X1 U334 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U335 ( .A(G92GAT), .B(G85GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(n430), .B(KEYINPUT46), .ZN(n431) );
  XNOR2_X1 U337 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U338 ( .A(n435), .B(KEYINPUT47), .ZN(n436) );
  XNOR2_X1 U339 ( .A(n437), .B(n436), .ZN(n444) );
  XNOR2_X1 U340 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n458) );
  XNOR2_X1 U341 ( .A(G92GAT), .B(KEYINPUT98), .ZN(n447) );
  XNOR2_X1 U342 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U343 ( .A(n426), .B(n425), .ZN(n428) );
  AND2_X1 U344 ( .A1(n466), .A2(n527), .ZN(n465) );
  XNOR2_X1 U345 ( .A(n451), .B(n294), .ZN(n452) );
  XNOR2_X1 U346 ( .A(n439), .B(n429), .ZN(n559) );
  XNOR2_X1 U347 ( .A(n453), .B(n452), .ZN(n457) );
  INV_X1 U348 ( .A(G218GAT), .ZN(n462) );
  XNOR2_X1 U349 ( .A(n310), .B(n292), .ZN(n567) );
  XNOR2_X1 U350 ( .A(n462), .B(KEYINPUT62), .ZN(n463) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n491) );
  XNOR2_X1 U352 ( .A(n481), .B(G29GAT), .ZN(n482) );
  XNOR2_X1 U353 ( .A(n464), .B(n463), .ZN(G1355GAT) );
  XNOR2_X1 U354 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U355 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U357 ( .A(n295), .B(n296), .ZN(n410) );
  NAND2_X1 U358 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U359 ( .A(n293), .B(n297), .ZN(n302) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U361 ( .A(n298), .B(G218GAT), .ZN(n448) );
  XOR2_X1 U362 ( .A(KEYINPUT74), .B(n448), .Z(n300) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n347) );
  XNOR2_X1 U364 ( .A(G134GAT), .B(n347), .ZN(n299) );
  XNOR2_X1 U365 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U366 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n304) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U369 ( .A(KEYINPUT7), .B(n305), .ZN(n408) );
  INV_X1 U370 ( .A(n408), .ZN(n309) );
  XOR2_X1 U371 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n307) );
  XNOR2_X1 U372 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U374 ( .A(n567), .B(KEYINPUT75), .ZN(n549) );
  XNOR2_X1 U375 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n353) );
  XOR2_X1 U376 ( .A(G176GAT), .B(G190GAT), .Z(n312) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(G99GAT), .ZN(n311) );
  XNOR2_X1 U378 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U379 ( .A(KEYINPUT65), .B(KEYINPUT85), .Z(n314) );
  XNOR2_X1 U380 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n313) );
  XNOR2_X1 U381 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U382 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U383 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n318) );
  NAND2_X1 U384 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U385 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U386 ( .A(KEYINPUT20), .B(n319), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G127GAT), .Z(n379) );
  XOR2_X1 U389 ( .A(n322), .B(n379), .Z(n325) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(G134GAT), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n323), .B(KEYINPUT0), .ZN(n363) );
  XOR2_X1 U392 ( .A(G120GAT), .B(G71GAT), .Z(n416) );
  XNOR2_X1 U393 ( .A(n363), .B(n416), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n325), .B(n324), .ZN(n330) );
  XOR2_X1 U395 ( .A(KEYINPUT83), .B(G183GAT), .Z(n327) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n326) );
  XNOR2_X1 U397 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U398 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n328) );
  XOR2_X1 U399 ( .A(n329), .B(n328), .Z(n455) );
  XNOR2_X1 U400 ( .A(n330), .B(n455), .ZN(n541) );
  INV_X1 U401 ( .A(n541), .ZN(n531) );
  XOR2_X1 U402 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n332) );
  XNOR2_X1 U403 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n331) );
  XNOR2_X1 U404 ( .A(n332), .B(n331), .ZN(n338) );
  XOR2_X1 U405 ( .A(G211GAT), .B(KEYINPUT21), .Z(n334) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n333) );
  XNOR2_X1 U407 ( .A(n334), .B(n333), .ZN(n454) );
  XOR2_X1 U408 ( .A(KEYINPUT88), .B(n454), .Z(n336) );
  NAND2_X1 U409 ( .A1(G228GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U410 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n351) );
  XOR2_X1 U412 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n340) );
  XNOR2_X1 U413 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n339) );
  XNOR2_X1 U414 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U415 ( .A(n341), .B(G106GAT), .Z(n343) );
  XOR2_X1 U416 ( .A(G148GAT), .B(G78GAT), .Z(n423) );
  XNOR2_X1 U417 ( .A(n423), .B(G218GAT), .ZN(n342) );
  XNOR2_X1 U418 ( .A(n343), .B(n342), .ZN(n346) );
  XOR2_X1 U419 ( .A(G155GAT), .B(KEYINPUT2), .Z(n345) );
  XNOR2_X1 U420 ( .A(KEYINPUT3), .B(KEYINPUT90), .ZN(n344) );
  XNOR2_X1 U421 ( .A(n345), .B(n344), .ZN(n362) );
  XOR2_X1 U422 ( .A(n346), .B(n362), .Z(n349) );
  XOR2_X1 U423 ( .A(G141GAT), .B(G22GAT), .Z(n399) );
  XNOR2_X1 U424 ( .A(n399), .B(n347), .ZN(n348) );
  XNOR2_X1 U425 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U426 ( .A(n351), .B(n350), .ZN(n484) );
  NOR2_X1 U427 ( .A1(n531), .A2(n484), .ZN(n352) );
  XNOR2_X1 U428 ( .A(n353), .B(n352), .ZN(n554) );
  XOR2_X1 U429 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n355) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n354) );
  XNOR2_X1 U431 ( .A(n355), .B(n354), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n357) );
  XNOR2_X1 U433 ( .A(G127GAT), .B(KEYINPUT6), .ZN(n356) );
  XNOR2_X1 U434 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U435 ( .A(G57GAT), .B(KEYINPUT95), .Z(n359) );
  XNOR2_X1 U436 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n358) );
  XNOR2_X1 U437 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U438 ( .A(n361), .B(n360), .Z(n365) );
  XNOR2_X1 U439 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U440 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n367), .B(n366), .ZN(n375) );
  NAND2_X1 U442 ( .A1(G225GAT), .A2(G233GAT), .ZN(n373) );
  XOR2_X1 U443 ( .A(G148GAT), .B(G162GAT), .Z(n369) );
  XNOR2_X1 U444 ( .A(G141GAT), .B(G120GAT), .ZN(n368) );
  XNOR2_X1 U445 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U446 ( .A(G29GAT), .B(G85GAT), .Z(n370) );
  XNOR2_X1 U447 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U448 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n527) );
  XOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT76), .Z(n450) );
  XOR2_X1 U451 ( .A(n450), .B(G78GAT), .Z(n377) );
  XOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT69), .Z(n398) );
  XNOR2_X1 U453 ( .A(n398), .B(G155GAT), .ZN(n376) );
  XNOR2_X1 U454 ( .A(n377), .B(n376), .ZN(n383) );
  XNOR2_X1 U455 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n378) );
  XNOR2_X1 U456 ( .A(n378), .B(KEYINPUT13), .ZN(n422) );
  XOR2_X1 U457 ( .A(n422), .B(n379), .Z(n381) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U459 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U460 ( .A(n383), .B(n382), .Z(n385) );
  XNOR2_X1 U461 ( .A(G22GAT), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n385), .B(n384), .ZN(n393) );
  XOR2_X1 U463 ( .A(KEYINPUT78), .B(G64GAT), .Z(n387) );
  XNOR2_X1 U464 ( .A(G183GAT), .B(G71GAT), .ZN(n386) );
  XNOR2_X1 U465 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U466 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n389) );
  XNOR2_X1 U467 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U468 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U469 ( .A(n391), .B(n390), .Z(n392) );
  XNOR2_X1 U470 ( .A(n393), .B(n392), .ZN(n587) );
  XOR2_X1 U471 ( .A(G15GAT), .B(G113GAT), .Z(n395) );
  XNOR2_X1 U472 ( .A(G169GAT), .B(G197GAT), .ZN(n394) );
  XNOR2_X1 U473 ( .A(n395), .B(n394), .ZN(n407) );
  XOR2_X1 U474 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n397) );
  XNOR2_X1 U475 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n396) );
  XNOR2_X1 U476 ( .A(n397), .B(n396), .ZN(n403) );
  XOR2_X1 U477 ( .A(G50GAT), .B(G36GAT), .Z(n401) );
  XNOR2_X1 U478 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U479 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U480 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U481 ( .A1(G229GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U482 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U483 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U484 ( .A(n409), .B(n408), .Z(n515) );
  INV_X1 U485 ( .A(n515), .ZN(n578) );
  XNOR2_X1 U486 ( .A(n410), .B(KEYINPUT71), .ZN(n413) );
  INV_X1 U487 ( .A(n413), .ZN(n412) );
  INV_X1 U488 ( .A(KEYINPUT33), .ZN(n411) );
  NAND2_X1 U489 ( .A1(n412), .A2(n411), .ZN(n415) );
  NAND2_X1 U490 ( .A1(n413), .A2(KEYINPUT33), .ZN(n414) );
  NAND2_X1 U491 ( .A1(n415), .A2(n414), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n416), .B(KEYINPUT32), .ZN(n417) );
  XNOR2_X1 U493 ( .A(n417), .B(KEYINPUT31), .ZN(n418) );
  XNOR2_X1 U494 ( .A(n419), .B(n418), .ZN(n426) );
  XOR2_X1 U495 ( .A(G64GAT), .B(KEYINPUT72), .Z(n421) );
  XNOR2_X1 U496 ( .A(G176GAT), .B(G204GAT), .ZN(n420) );
  XNOR2_X1 U497 ( .A(n421), .B(n420), .ZN(n451) );
  XNOR2_X1 U498 ( .A(n451), .B(n422), .ZN(n424) );
  NAND2_X1 U499 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U500 ( .A(n428), .B(n427), .ZN(n439) );
  AND2_X1 U501 ( .A1(n578), .A2(n559), .ZN(n432) );
  INV_X1 U502 ( .A(KEYINPUT111), .ZN(n430) );
  NOR2_X1 U503 ( .A1(n587), .A2(n433), .ZN(n434) );
  NAND2_X1 U504 ( .A1(n434), .A2(n567), .ZN(n437) );
  XOR2_X1 U505 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n435) );
  INV_X1 U506 ( .A(n587), .ZN(n493) );
  NOR2_X1 U507 ( .A1(n493), .A2(n476), .ZN(n438) );
  XNOR2_X1 U508 ( .A(KEYINPUT45), .B(n438), .ZN(n440) );
  NAND2_X1 U509 ( .A1(n440), .A2(n439), .ZN(n441) );
  NOR2_X1 U510 ( .A1(n578), .A2(n441), .ZN(n442) );
  XNOR2_X1 U511 ( .A(KEYINPUT114), .B(n442), .ZN(n443) );
  NOR2_X1 U512 ( .A1(n444), .A2(n443), .ZN(n446) );
  INV_X1 U513 ( .A(KEYINPUT48), .ZN(n445) );
  XNOR2_X1 U514 ( .A(n446), .B(n445), .ZN(n538) );
  XOR2_X1 U515 ( .A(n450), .B(n449), .Z(n453) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(n529) );
  NAND2_X1 U518 ( .A1(n538), .A2(n529), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n554), .A2(n485), .ZN(n461) );
  INV_X1 U520 ( .A(n586), .ZN(n583) );
  NOR2_X1 U521 ( .A1(n476), .A2(n583), .ZN(n464) );
  XOR2_X1 U522 ( .A(n484), .B(KEYINPUT28), .Z(n533) );
  XNOR2_X1 U523 ( .A(n529), .B(KEYINPUT27), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n533), .A2(n556), .ZN(n539) );
  NAND2_X1 U525 ( .A1(n539), .A2(n541), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n466), .A2(n554), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n531), .A2(n529), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n484), .A2(n467), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NAND2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n472) );
  INV_X1 U531 ( .A(n527), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT101), .ZN(n497) );
  NOR2_X1 U535 ( .A1(n497), .A2(n476), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n477), .A2(n493), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT37), .B(n478), .Z(n526) );
  NAND2_X1 U538 ( .A1(n439), .A2(n578), .ZN(n498) );
  NOR2_X1 U539 ( .A1(n526), .A2(n498), .ZN(n479) );
  XOR2_X1 U540 ( .A(KEYINPUT105), .B(n479), .Z(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT38), .B(n480), .ZN(n513) );
  NAND2_X1 U542 ( .A1(n527), .A2(n513), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n481) );
  INV_X1 U544 ( .A(KEYINPUT122), .ZN(n490) );
  NAND2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n488), .A2(n531), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n576) );
  NAND2_X1 U550 ( .A1(n576), .A2(n549), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n495) );
  OR2_X1 U552 ( .A1(n549), .A2(n493), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  OR2_X1 U554 ( .A1(n497), .A2(n496), .ZN(n516) );
  NOR2_X1 U555 ( .A1(n498), .A2(n516), .ZN(n499) );
  XNOR2_X1 U556 ( .A(KEYINPUT102), .B(n499), .ZN(n507) );
  NAND2_X1 U557 ( .A1(n507), .A2(n527), .ZN(n502) );
  XOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT34), .Z(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT103), .B(n500), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n507), .A2(n529), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U564 ( .A1(n531), .A2(n507), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n533), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(G36GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U570 ( .A1(n529), .A2(n513), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n531), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n533), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U578 ( .A(n559), .B(KEYINPUT108), .ZN(n573) );
  NAND2_X1 U579 ( .A1(n515), .A2(n573), .ZN(n525) );
  NOR2_X1 U580 ( .A1(n516), .A2(n525), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n527), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n529), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n531), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n536) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n537), .Z(G1339GAT) );
  XOR2_X1 U602 ( .A(G113GAT), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U603 ( .A1(n538), .A2(n539), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n550), .A2(n578), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U608 ( .A1(n550), .A2(n573), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U611 ( .A1(n550), .A2(n587), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  NAND2_X1 U618 ( .A1(n538), .A2(n554), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n578), .A2(n565), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT118), .ZN(n558) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n558), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  NAND2_X1 U624 ( .A1(n565), .A2(n559), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT119), .Z(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n587), .A2(n565), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U630 ( .A(n565), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n576), .A2(n578), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(n572), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n576), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n586), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  OR2_X1 U649 ( .A1(n583), .A2(n439), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
endmodule

