//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT73), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT75), .ZN(new_n202));
  OR3_X1    g016(.A1(new_n195), .A2(KEYINPUT75), .A3(G125), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G119), .B(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT74), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT24), .B(G110), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G128), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n212), .A2(G128), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(new_n215), .C1(new_n216), .C2(KEYINPUT23), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT76), .B(G110), .Z(new_n218));
  OR2_X1    g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI211_X1 g033(.A(new_n200), .B(new_n207), .C1(new_n211), .C2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n204), .A2(new_n201), .A3(new_n206), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(G110), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n209), .B2(new_n210), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n194), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n211), .A2(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n204), .A2(new_n206), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  INV_X1    g043(.A(new_n200), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI221_X1 g045(.A(new_n223), .B1(new_n209), .B2(new_n210), .C1(new_n221), .C2(new_n207), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n193), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n233), .A3(new_n188), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n189), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n189), .A2(G902), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n239), .A3(new_n233), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G134), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n243), .A2(G137), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n255));
  OAI211_X1 g069(.A(KEYINPUT67), .B(new_n246), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT68), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n248), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n250), .A2(new_n249), .A3(new_n251), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT67), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n260), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(KEYINPUT68), .A3(G131), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n201), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G146), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT65), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n272), .ZN(new_n278));
  NOR2_X1   g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n275), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n269), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n265), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n278), .A2(new_n285), .A3(G128), .ZN(new_n286));
  INV_X1    g100(.A(new_n244), .ZN(new_n287));
  OAI21_X1  g101(.A(G131), .B1(new_n287), .B2(new_n251), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n270), .B(new_n272), .C1(KEYINPUT1), .C2(new_n214), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n283), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n284), .B1(new_n283), .B2(new_n290), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT2), .B(G113), .Z(new_n297));
  XNOR2_X1  g111(.A(G116), .B(G119), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n283), .A2(new_n290), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n282), .A2(KEYINPUT30), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n296), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n301), .B(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(KEYINPUT71), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n304), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n304), .A2(new_n314), .A3(KEYINPUT31), .A4(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n306), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n282), .A2(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT28), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n311), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT32), .ZN(new_n330));
  NOR2_X1   g144(.A1(G472), .A2(G902), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n318), .A2(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n333));
  INV_X1    g147(.A(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT32), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n304), .A2(new_n306), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n311), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n326), .B2(new_n327), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n188), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n282), .A2(new_n302), .ZN(new_n343));
  INV_X1    g157(.A(new_n305), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n306), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(KEYINPUT72), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(KEYINPUT28), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n325), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(new_n340), .A3(new_n327), .ZN(new_n351));
  OAI21_X1  g165(.A(G472), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n242), .B1(new_n336), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n298), .A2(KEYINPUT5), .ZN(new_n354));
  INV_X1    g168(.A(G116), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n355), .A2(KEYINPUT5), .A3(G119), .ZN(new_n356));
  INV_X1    g170(.A(G113), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n300), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(new_n361), .B2(G107), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G104), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(G107), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n361), .A2(G107), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n364), .A2(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(G101), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT89), .B1(new_n360), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n354), .A2(new_n358), .B1(new_n297), .B2(new_n298), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n360), .A2(new_n372), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT8), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n374), .A2(new_n375), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n362), .A2(new_n365), .A3(new_n367), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G101), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n301), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT81), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n366), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n384), .A2(KEYINPUT82), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT82), .B1(new_n384), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n380), .B(new_n383), .C1(new_n387), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n275), .A2(new_n277), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n278), .A2(new_n280), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(G125), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT88), .B1(new_n281), .B2(new_n197), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n286), .A2(new_n289), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n197), .ZN(new_n403));
  INV_X1    g217(.A(G224), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT7), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n401), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n382), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(KEYINPUT90), .A3(new_n197), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n400), .A2(new_n401), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n406), .B2(new_n405), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n405), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n383), .B1(new_n387), .B2(new_n395), .ZN(new_n418));
  INV_X1    g232(.A(new_n380), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT91), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n415), .A2(new_n426), .A3(new_n424), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  OAI21_X1  g248(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT78), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n188), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n268), .A2(new_n269), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n386), .A2(new_n281), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT83), .B1(new_n441), .B2(new_n395), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n384), .A2(new_n392), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n384), .A2(new_n392), .A3(KEYINPUT82), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n281), .A4(new_n386), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n402), .A2(new_n372), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n402), .B2(new_n372), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n442), .A2(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n440), .B1(new_n455), .B2(KEYINPUT85), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n449), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n454), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n457), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT86), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n458), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(KEYINPUT85), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n440), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n439), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT79), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT80), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n191), .A2(G227), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n402), .B(new_n372), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n268), .A2(new_n269), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n478), .A2(new_n479), .B1(new_n455), .B2(new_n439), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(KEYINPUT12), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(KEYINPUT87), .A3(new_n473), .A4(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n268), .A2(new_n479), .A3(new_n269), .A4(new_n476), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n467), .A2(new_n473), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g301(.A(G469), .B(new_n438), .C1(new_n475), .C2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n460), .A2(new_n466), .A3(new_n467), .A4(new_n473), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n474), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(G469), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G469), .A2(G902), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n433), .B(new_n437), .C1(new_n488), .C2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n361), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  INV_X1    g313(.A(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n191), .A3(G214), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n271), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n258), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n258), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n503), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G131), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT93), .A3(new_n504), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n229), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n202), .A2(new_n203), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT92), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(KEYINPUT94), .A3(KEYINPUT19), .A4(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n202), .A2(KEYINPUT92), .A3(new_n203), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT92), .B1(new_n202), .B2(new_n203), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT19), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n199), .B2(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n516), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n511), .B1(new_n523), .B2(new_n201), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n514), .A2(G146), .A3(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n230), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n508), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n498), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT95), .B1(new_n222), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n204), .A2(new_n201), .A3(new_n206), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n229), .A2(KEYINPUT95), .A3(new_n534), .A4(new_n532), .ZN(new_n535));
  OR3_X1    g349(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n529), .B(new_n497), .C1(new_n533), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n540));
  OR3_X1    g354(.A1(new_n540), .A2(G475), .A3(G902), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(G475), .B2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(KEYINPUT98), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(KEYINPUT98), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n539), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n531), .A2(KEYINPUT96), .A3(new_n538), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n543), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n553), .B2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(G475), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n529), .B1(new_n533), .B2(new_n537), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n498), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G902), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n558), .A3(new_n538), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  AOI211_X1 g378(.A(G953), .B(new_n564), .C1(G234), .C2(G237), .ZN(new_n565));
  AOI211_X1 g379(.A(new_n191), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT21), .B(G898), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n434), .A2(new_n187), .A3(G953), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n355), .A2(G122), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n355), .A2(G122), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n573), .B2(KEYINPUT14), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n575), .B2(new_n574), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(G107), .ZN(new_n578));
  INV_X1    g392(.A(new_n571), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n579), .A2(G107), .A3(new_n573), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n271), .A2(G128), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n214), .A2(G143), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n243), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n243), .B1(new_n582), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n589), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n582), .A2(new_n588), .A3(new_n589), .ZN(new_n593));
  OAI21_X1  g407(.A(G134), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G107), .B1(new_n579), .B2(new_n573), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n581), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n584), .ZN(new_n599));
  OAI221_X1 g413(.A(new_n570), .B1(new_n578), .B2(new_n587), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n570), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n594), .A2(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(KEYINPUT101), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n578), .A2(new_n587), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n188), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n563), .A2(new_n569), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n495), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n353), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  AOI21_X1  g430(.A(new_n438), .B1(new_n320), .B2(new_n328), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(new_n334), .B2(new_n333), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n475), .A2(new_n487), .ZN(new_n621));
  INV_X1    g435(.A(G469), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n188), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n492), .A2(new_n493), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n436), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n241), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n426), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n425), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n429), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n415), .A2(new_n424), .A3(KEYINPUT103), .A4(new_n426), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n431), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n548), .ZN(new_n636));
  INV_X1    g450(.A(new_n562), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT33), .B1(new_n570), .B2(KEYINPUT104), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n607), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n600), .A2(new_n606), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n640), .A2(G478), .A3(new_n188), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n608), .A2(new_n609), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n634), .A2(new_n638), .A3(new_n569), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n626), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NOR2_X1   g463(.A1(new_n612), .A2(new_n562), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n553), .B(KEYINPUT20), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n634), .A2(new_n650), .A3(new_n569), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n626), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n495), .A2(new_n619), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n231), .A2(new_n232), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n239), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n238), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n613), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  NAND2_X1  g479(.A1(new_n238), .A2(new_n660), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n630), .A2(new_n632), .A3(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n436), .B(new_n667), .C1(new_n623), .C2(new_n624), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n352), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n565), .ZN(new_n673));
  INV_X1    g487(.A(new_n566), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(G900), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n650), .A2(new_n651), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XNOR2_X1  g493(.A(new_n675), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n625), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT40), .Z(new_n682));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n347), .A2(new_n327), .A3(new_n348), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n316), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n336), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n611), .B1(new_n554), .B2(new_n562), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n430), .B(KEYINPUT38), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n661), .A2(new_n431), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n684), .A2(new_n685), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  OAI211_X1 g510(.A(new_n645), .B(new_n675), .C1(new_n554), .C2(new_n562), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n672), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(G146), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G48));
  NAND2_X1  g515(.A1(new_n482), .A2(new_n486), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n468), .B2(new_n474), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(new_n438), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n623), .A3(new_n435), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n646), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n353), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NOR2_X1   g523(.A1(new_n652), .A2(new_n705), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n353), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NOR2_X1   g526(.A1(new_n705), .A2(new_n633), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n671), .A3(new_n662), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  XNOR2_X1  g529(.A(KEYINPUT109), .B(G472), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n333), .B2(new_n438), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n350), .A2(new_n327), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n320), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n331), .B(KEYINPUT108), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n721), .A3(new_n241), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n717), .A2(new_n721), .A3(KEYINPUT110), .A4(new_n241), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n704), .A2(new_n569), .A3(new_n623), .A4(new_n435), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n634), .A2(new_n638), .A3(KEYINPUT111), .A4(new_n611), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n691), .B2(new_n633), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  AND3_X1   g547(.A1(new_n717), .A2(new_n721), .A3(new_n666), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n713), .A2(new_n698), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND4_X1  g550(.A1(new_n638), .A2(KEYINPUT106), .A3(new_n645), .A4(new_n675), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n697), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT114), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n737), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n430), .A2(new_n431), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n493), .B(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n492), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n435), .B1(new_n488), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n435), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n492), .A2(new_n744), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n623), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n353), .A2(new_n742), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n740), .A2(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n743), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n751), .B2(KEYINPUT113), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n746), .A2(new_n747), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n754), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n353), .A3(new_n742), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n258), .ZN(G33));
  NAND4_X1  g577(.A1(new_n353), .A2(new_n748), .A3(new_n677), .A4(new_n752), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT115), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NAND2_X1  g580(.A1(new_n563), .A2(new_n645), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT43), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n768), .A2(new_n620), .A3(new_n661), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n743), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n489), .B2(new_n491), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n622), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n491), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n744), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n623), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n435), .A3(new_n680), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n771), .B(new_n782), .C1(new_n770), .C2(new_n769), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n435), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(KEYINPUT47), .A3(new_n435), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n671), .A2(new_n241), .A3(new_n743), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n698), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NOR2_X1   g606(.A1(new_n768), .A2(new_n673), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n705), .A2(new_n743), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n734), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n242), .A2(new_n673), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n638), .A2(new_n645), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n690), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n692), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n431), .A3(new_n705), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n793), .A2(new_n726), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n793), .A2(new_n726), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n743), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n704), .A2(new_n623), .A3(new_n436), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT121), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n789), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n690), .A2(new_n794), .A3(new_n796), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n638), .A2(new_n645), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n564), .B(G953), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n713), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n793), .A2(new_n353), .A3(new_n794), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n821));
  OAI221_X1 g635(.A(new_n817), .B1(new_n818), .B2(new_n808), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n824));
  INV_X1    g638(.A(new_n799), .ZN(new_n825));
  INV_X1    g639(.A(new_n806), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT51), .B(new_n825), .C1(new_n826), .C2(new_n804), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n787), .A2(new_n788), .A3(new_n810), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n809), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n824), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n807), .A2(KEYINPUT122), .A3(KEYINPUT51), .A4(new_n829), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n823), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n823), .B2(new_n833), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n353), .A2(new_n614), .B1(new_n656), .B2(new_n662), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n563), .A2(new_n612), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n644), .B(new_n643), .C1(new_n554), .C2(new_n562), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n569), .A2(new_n839), .A3(new_n433), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n241), .A3(new_n620), .A4(new_n625), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n748), .A2(new_n698), .A3(new_n734), .A4(new_n752), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n612), .A2(new_n666), .A3(new_n675), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n637), .A2(new_n756), .A3(new_n844), .A4(new_n651), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n671), .A3(new_n625), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n838), .A2(new_n842), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n353), .B1(new_n706), .B2(new_n710), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n732), .A2(new_n714), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n671), .B(new_n668), .C1(new_n698), .C2(new_n677), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n728), .A2(new_n730), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n675), .B(KEYINPUT118), .Z(new_n853));
  NAND2_X1  g667(.A1(new_n661), .A2(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n749), .B(new_n854), .C1(new_n623), .C2(new_n750), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n689), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n735), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n851), .A2(new_n856), .A3(new_n735), .A4(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n755), .A2(new_n761), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n850), .A2(new_n861), .A3(new_n862), .A4(new_n765), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n764), .A2(KEYINPUT115), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n764), .A2(KEYINPUT115), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n762), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n861), .A4(new_n850), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(KEYINPUT120), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n868), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n864), .B2(new_n869), .ZN(new_n877));
  AND4_X1   g691(.A1(KEYINPUT117), .A2(new_n863), .A3(new_n868), .A4(new_n861), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n879), .B2(KEYINPUT54), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT119), .A4(new_n871), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n837), .B(new_n874), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n564), .A2(new_n191), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n767), .A2(new_n242), .A3(new_n432), .A4(new_n436), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT116), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n704), .A2(new_n623), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT49), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n800), .B1(new_n887), .B2(KEYINPUT49), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n886), .A2(new_n690), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n421), .A2(new_n423), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n417), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n870), .A2(new_n188), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n627), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n191), .A2(G952), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n897), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n895), .B2(new_n427), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(G51));
  XNOR2_X1  g716(.A(new_n870), .B(new_n871), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n744), .B(KEYINPUT57), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n621), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n774), .A3(new_n773), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n551), .A2(new_n552), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n899), .ZN(G60));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT59), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n903), .A2(new_n640), .A3(new_n642), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n899), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n640), .A2(new_n642), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT60), .Z(new_n924));
  NAND3_X1  g738(.A1(new_n864), .A2(new_n869), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n226), .A2(new_n233), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n899), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n864), .A2(new_n869), .A3(new_n659), .A4(new_n924), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(KEYINPUT61), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n932), .A2(KEYINPUT125), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT125), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(G66));
  NAND2_X1  g750(.A1(new_n838), .A2(new_n842), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n849), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n191), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n567), .B2(new_n404), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n892), .B1(G898), .B2(new_n191), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  NAND2_X1  g757(.A1(new_n296), .A2(new_n303), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n523), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n851), .A2(new_n735), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n695), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n839), .A2(new_n840), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n681), .A2(new_n743), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n353), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n948), .B2(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n783), .A2(new_n791), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n945), .B1(new_n955), .B2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n191), .A2(G900), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n353), .A2(new_n852), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n946), .B1(new_n782), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n867), .A2(new_n783), .A3(new_n791), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n960), .B2(new_n191), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g776(.A(new_n945), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n961), .B2(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n956), .B(new_n968), .C1(new_n962), .C2(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  NOR4_X1   g784(.A1(new_n949), .A2(new_n953), .A3(new_n938), .A4(new_n954), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT63), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n311), .B(new_n337), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n960), .A2(new_n938), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n327), .B(new_n338), .C1(new_n975), .C2(new_n973), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n917), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n339), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n978), .B2(new_n316), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n879), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(G57));
endmodule


