

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741;

  NOR2_X1 U364 ( .A1(n666), .A2(n663), .ZN(n695) );
  NOR2_X1 U365 ( .A1(n607), .A2(n468), .ZN(n429) );
  XNOR2_X1 U366 ( .A(n429), .B(n428), .ZN(n557) );
  XNOR2_X2 U367 ( .A(G101), .B(G110), .ZN(n415) );
  XNOR2_X2 U368 ( .A(n359), .B(G143), .ZN(n440) );
  XNOR2_X2 U369 ( .A(G128), .B(KEYINPUT65), .ZN(n359) );
  INV_X1 U370 ( .A(n523), .ZN(n371) );
  OR2_X2 U371 ( .A1(n523), .A2(n677), .ZN(n530) );
  NAND2_X1 U372 ( .A1(n406), .A2(n405), .ZN(n404) );
  AND2_X1 U373 ( .A1(n605), .A2(n346), .ZN(n405) );
  XNOR2_X1 U374 ( .A(n394), .B(n393), .ZN(n605) );
  AND2_X1 U375 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U376 ( .A1(n348), .A2(n385), .ZN(n378) );
  NOR2_X1 U377 ( .A1(n544), .A2(KEYINPUT44), .ZN(n545) );
  XNOR2_X1 U378 ( .A(n386), .B(KEYINPUT106), .ZN(n741) );
  NOR2_X1 U379 ( .A1(n541), .A2(n514), .ZN(n516) );
  NAND2_X1 U380 ( .A1(n517), .A2(n590), .ZN(n541) );
  INV_X2 U381 ( .A(G953), .ZN(n731) );
  XNOR2_X1 U382 ( .A(KEYINPUT100), .B(n343), .ZN(n535) );
  NAND2_X1 U383 ( .A1(n534), .A2(n555), .ZN(n343) );
  NAND2_X1 U384 ( .A1(n392), .A2(n389), .ZN(n388) );
  BUF_X1 U385 ( .A(n631), .Z(n344) );
  XNOR2_X1 U386 ( .A(n516), .B(n515), .ZN(n631) );
  AND2_X1 U387 ( .A1(n546), .A2(n616), .ZN(n345) );
  NOR2_X2 U388 ( .A1(n631), .A2(n617), .ZN(n546) );
  XNOR2_X2 U389 ( .A(n388), .B(n354), .ZN(n720) );
  OR2_X2 U390 ( .A1(n713), .A2(n356), .ZN(n628) );
  XNOR2_X1 U391 ( .A(n440), .B(KEYINPUT4), .ZN(n475) );
  OR2_X1 U392 ( .A1(n644), .A2(G902), .ZN(n496) );
  XNOR2_X1 U393 ( .A(n475), .B(n474), .ZN(n489) );
  XNOR2_X1 U394 ( .A(n397), .B(n513), .ZN(n674) );
  INV_X1 U395 ( .A(n695), .ZN(n387) );
  INV_X1 U396 ( .A(KEYINPUT69), .ZN(n391) );
  XNOR2_X1 U397 ( .A(n459), .B(n409), .ZN(n412) );
  XNOR2_X1 U398 ( .A(n410), .B(KEYINPUT17), .ZN(n411) );
  NAND2_X1 U399 ( .A1(n524), .A2(n369), .ZN(n368) );
  NAND2_X1 U400 ( .A1(n371), .A2(n370), .ZN(n369) );
  NOR2_X1 U401 ( .A1(n677), .A2(KEYINPUT33), .ZN(n370) );
  XNOR2_X1 U402 ( .A(KEYINPUT16), .B(G122), .ZN(n421) );
  XNOR2_X1 U403 ( .A(n489), .B(n358), .ZN(n357) );
  INV_X1 U404 ( .A(n713), .ZN(n362) );
  NAND2_X1 U405 ( .A1(n557), .A2(n690), .ZN(n401) );
  NAND2_X1 U406 ( .A1(n570), .A2(n569), .ZN(n398) );
  NOR2_X1 U407 ( .A1(n587), .A2(n566), .ZN(n567) );
  XNOR2_X1 U408 ( .A(n467), .B(n466), .ZN(n538) );
  XNOR2_X1 U409 ( .A(n465), .B(n464), .ZN(n466) );
  INV_X1 U410 ( .A(KEYINPUT91), .ZN(n379) );
  XOR2_X1 U411 ( .A(G104), .B(G113), .Z(n452) );
  NAND2_X1 U412 ( .A1(n565), .A2(n674), .ZN(n587) );
  AND2_X1 U413 ( .A1(n561), .A2(n471), .ZN(n472) );
  INV_X1 U414 ( .A(G137), .ZN(n479) );
  XNOR2_X1 U415 ( .A(G128), .B(G119), .ZN(n501) );
  XNOR2_X1 U416 ( .A(n400), .B(n399), .ZN(n498) );
  INV_X1 U417 ( .A(KEYINPUT8), .ZN(n399) );
  NAND2_X1 U418 ( .A1(n731), .A2(G234), .ZN(n400) );
  XNOR2_X1 U419 ( .A(G134), .B(G116), .ZN(n445) );
  XNOR2_X1 U420 ( .A(n412), .B(n411), .ZN(n413) );
  INV_X1 U421 ( .A(KEYINPUT48), .ZN(n393) );
  NAND2_X1 U422 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U423 ( .A1(n530), .A2(KEYINPUT33), .ZN(n365) );
  NAND2_X1 U424 ( .A1(n590), .A2(n372), .ZN(n367) );
  INV_X1 U425 ( .A(G472), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n357), .B(n347), .ZN(n644) );
  NAND2_X1 U427 ( .A1(n362), .A2(n360), .ZN(n611) );
  INV_X1 U428 ( .A(G210), .ZN(n361) );
  NOR2_X1 U429 ( .A1(n398), .A2(n580), .ZN(n661) );
  NOR2_X1 U430 ( .A1(n540), .A2(n539), .ZN(n663) );
  NAND2_X1 U431 ( .A1(n373), .A2(n351), .ZN(n386) );
  INV_X1 U432 ( .A(n543), .ZN(n373) );
  AND2_X1 U433 ( .A1(n604), .A2(KEYINPUT2), .ZN(n346) );
  XOR2_X1 U434 ( .A(n494), .B(n493), .Z(n347) );
  AND2_X1 U435 ( .A1(n384), .A2(n379), .ZN(n348) );
  OR2_X1 U436 ( .A1(n665), .A2(n652), .ZN(n349) );
  AND2_X1 U437 ( .A1(n374), .A2(KEYINPUT91), .ZN(n350) );
  AND2_X1 U438 ( .A1(n523), .A2(n542), .ZN(n351) );
  NOR2_X1 U439 ( .A1(n707), .A2(n398), .ZN(n352) );
  NAND2_X1 U440 ( .A1(n366), .A2(n365), .ZN(n699) );
  XOR2_X1 U441 ( .A(KEYINPUT22), .B(KEYINPUT76), .Z(n353) );
  INV_X1 U442 ( .A(KEYINPUT33), .ZN(n372) );
  XOR2_X1 U443 ( .A(n547), .B(KEYINPUT64), .Z(n354) );
  XOR2_X1 U444 ( .A(KEYINPUT46), .B(KEYINPUT89), .Z(n355) );
  INV_X1 U445 ( .A(KEYINPUT2), .ZN(n408) );
  OR2_X1 U446 ( .A1(n606), .A2(n364), .ZN(n356) );
  INV_X1 U447 ( .A(G475), .ZN(n464) );
  XNOR2_X1 U448 ( .A(n357), .B(n729), .ZN(n733) );
  INV_X1 U449 ( .A(n503), .ZN(n358) );
  NAND2_X1 U450 ( .A1(n362), .A2(n363), .ZN(n620) );
  NOR2_X1 U451 ( .A1(n713), .A2(n606), .ZN(n642) );
  NOR2_X1 U452 ( .A1(n606), .A2(n361), .ZN(n360) );
  NOR2_X1 U453 ( .A1(n606), .A2(n464), .ZN(n363) );
  NAND2_X1 U454 ( .A1(n529), .A2(KEYINPUT44), .ZN(n385) );
  NAND2_X1 U455 ( .A1(n376), .A2(n350), .ZN(n381) );
  NAND2_X1 U456 ( .A1(n384), .A2(n375), .ZN(n374) );
  INV_X1 U457 ( .A(KEYINPUT44), .ZN(n375) );
  NAND2_X1 U458 ( .A1(n345), .A2(n384), .ZN(n376) );
  NAND2_X1 U459 ( .A1(n380), .A2(n377), .ZN(n392) );
  NAND2_X1 U460 ( .A1(n378), .A2(n741), .ZN(n377) );
  NAND2_X1 U461 ( .A1(n383), .A2(KEYINPUT91), .ZN(n382) );
  INV_X1 U462 ( .A(n741), .ZN(n383) );
  NAND2_X1 U463 ( .A1(n349), .A2(n387), .ZN(n384) );
  NAND2_X1 U464 ( .A1(n390), .A2(n546), .ZN(n389) );
  XNOR2_X1 U465 ( .A(n545), .B(n391), .ZN(n390) );
  NAND2_X1 U466 ( .A1(n605), .A2(n604), .ZN(n730) );
  NAND2_X1 U467 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n595), .B(KEYINPUT72), .ZN(n395) );
  XNOR2_X1 U469 ( .A(n571), .B(n355), .ZN(n396) );
  NAND2_X1 U470 ( .A1(n632), .A2(n509), .ZN(n397) );
  XNOR2_X2 U471 ( .A(n586), .B(KEYINPUT19), .ZN(n579) );
  XNOR2_X2 U472 ( .A(n401), .B(KEYINPUT93), .ZN(n586) );
  AND2_X2 U473 ( .A1(n403), .A2(n402), .ZN(n407) );
  NAND2_X1 U474 ( .A1(n730), .A2(n408), .ZN(n402) );
  NAND2_X1 U475 ( .A1(n720), .A2(n408), .ZN(n403) );
  NAND2_X2 U476 ( .A1(n407), .A2(n404), .ZN(n713) );
  INV_X1 U477 ( .A(n720), .ZN(n406) );
  XNOR2_X2 U478 ( .A(KEYINPUT3), .B(G119), .ZN(n419) );
  INV_X1 U479 ( .A(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U480 ( .A(G113), .B(G116), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U482 ( .A(G104), .B(G107), .ZN(n414) );
  NOR2_X1 U483 ( .A1(G953), .A2(G237), .ZN(n476) );
  INV_X1 U484 ( .A(n522), .ZN(n471) );
  XNOR2_X1 U485 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U486 ( .A(KEYINPUT99), .ZN(n532) );
  BUF_X1 U487 ( .A(n557), .Z(n600) );
  XOR2_X2 U488 ( .A(G146), .B(G125), .Z(n459) );
  NAND2_X1 U489 ( .A1(G224), .A2(n731), .ZN(n410) );
  XNOR2_X1 U490 ( .A(n475), .B(n413), .ZN(n423) );
  INV_X1 U491 ( .A(n414), .ZN(n416) );
  XNOR2_X2 U492 ( .A(n416), .B(n415), .ZN(n715) );
  XNOR2_X1 U493 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n417) );
  XNOR2_X2 U494 ( .A(n715), .B(n417), .ZN(n494) );
  INV_X1 U495 ( .A(n418), .ZN(n420) );
  XNOR2_X2 U496 ( .A(n420), .B(n419), .ZN(n484) );
  XNOR2_X2 U497 ( .A(n484), .B(n421), .ZN(n716) );
  XNOR2_X1 U498 ( .A(n494), .B(n716), .ZN(n422) );
  XNOR2_X1 U499 ( .A(n422), .B(n423), .ZN(n607) );
  INV_X1 U500 ( .A(KEYINPUT15), .ZN(n424) );
  XNOR2_X1 U501 ( .A(n424), .B(G902), .ZN(n468) );
  XOR2_X1 U502 ( .A(KEYINPUT95), .B(KEYINPUT84), .Z(n427) );
  NOR2_X1 U503 ( .A1(G237), .A2(G902), .ZN(n425) );
  XOR2_X1 U504 ( .A(KEYINPUT78), .B(n425), .Z(n430) );
  NAND2_X1 U505 ( .A1(n430), .A2(G210), .ZN(n426) );
  XNOR2_X1 U506 ( .A(n427), .B(n426), .ZN(n428) );
  NAND2_X1 U507 ( .A1(n430), .A2(G214), .ZN(n690) );
  XOR2_X1 U508 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n432) );
  NAND2_X1 U509 ( .A1(G234), .A2(G237), .ZN(n431) );
  XNOR2_X1 U510 ( .A(n432), .B(n431), .ZN(n433) );
  NAND2_X1 U511 ( .A1(G952), .A2(n433), .ZN(n706) );
  NOR2_X1 U512 ( .A1(G953), .A2(n706), .ZN(n552) );
  NAND2_X1 U513 ( .A1(G902), .A2(n433), .ZN(n548) );
  INV_X1 U514 ( .A(n548), .ZN(n434) );
  NOR2_X1 U515 ( .A1(G898), .A2(n731), .ZN(n718) );
  NAND2_X1 U516 ( .A1(n434), .A2(n718), .ZN(n435) );
  XOR2_X1 U517 ( .A(KEYINPUT96), .B(n435), .Z(n436) );
  NOR2_X1 U518 ( .A1(n552), .A2(n436), .ZN(n437) );
  NOR2_X2 U519 ( .A1(n579), .A2(n437), .ZN(n439) );
  XNOR2_X1 U520 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n438) );
  XNOR2_X2 U521 ( .A(n439), .B(n438), .ZN(n534) );
  NAND2_X1 U522 ( .A1(n498), .A2(G217), .ZN(n441) );
  XNOR2_X1 U523 ( .A(n441), .B(n440), .ZN(n448) );
  XOR2_X1 U524 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n443) );
  XNOR2_X1 U525 ( .A(G107), .B(G122), .ZN(n442) );
  XNOR2_X1 U526 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U527 ( .A(n444), .B(KEYINPUT102), .Z(n446) );
  XNOR2_X1 U528 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U529 ( .A(n448), .B(n447), .ZN(n638) );
  INV_X1 U530 ( .A(G902), .ZN(n509) );
  NAND2_X1 U531 ( .A1(n638), .A2(n509), .ZN(n450) );
  XOR2_X1 U532 ( .A(KEYINPUT103), .B(G478), .Z(n449) );
  XNOR2_X1 U533 ( .A(n450), .B(n449), .ZN(n539) );
  XNOR2_X1 U534 ( .A(G143), .B(G131), .ZN(n451) );
  XNOR2_X1 U535 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n454) );
  XNOR2_X1 U537 ( .A(G122), .B(KEYINPUT12), .ZN(n453) );
  XNOR2_X1 U538 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U539 ( .A(n456), .B(n455), .Z(n458) );
  NAND2_X1 U540 ( .A1(G214), .A2(n476), .ZN(n457) );
  XNOR2_X1 U541 ( .A(n458), .B(n457), .ZN(n463) );
  XNOR2_X1 U542 ( .A(n459), .B(G140), .ZN(n461) );
  INV_X1 U543 ( .A(KEYINPUT10), .ZN(n460) );
  XNOR2_X1 U544 ( .A(n461), .B(n460), .ZN(n729) );
  INV_X1 U545 ( .A(n729), .ZN(n462) );
  XNOR2_X1 U546 ( .A(n463), .B(n462), .ZN(n618) );
  NOR2_X1 U547 ( .A1(G902), .A2(n618), .ZN(n467) );
  INV_X1 U548 ( .A(KEYINPUT13), .ZN(n465) );
  NOR2_X1 U549 ( .A1(n539), .A2(n538), .ZN(n561) );
  INV_X1 U550 ( .A(n468), .ZN(n606) );
  NAND2_X1 U551 ( .A1(G234), .A2(n606), .ZN(n469) );
  XNOR2_X1 U552 ( .A(KEYINPUT20), .B(n469), .ZN(n510) );
  NAND2_X1 U553 ( .A1(n510), .A2(G221), .ZN(n470) );
  XNOR2_X1 U554 ( .A(n470), .B(KEYINPUT21), .ZN(n673) );
  XNOR2_X1 U555 ( .A(n673), .B(KEYINPUT98), .ZN(n522) );
  NAND2_X1 U556 ( .A1(n534), .A2(n472), .ZN(n473) );
  XNOR2_X2 U557 ( .A(n473), .B(n353), .ZN(n517) );
  XNOR2_X1 U558 ( .A(G134), .B(G131), .ZN(n474) );
  XOR2_X1 U559 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n478) );
  NAND2_X1 U560 ( .A1(n476), .A2(G210), .ZN(n477) );
  XNOR2_X1 U561 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U562 ( .A(G101), .B(G146), .ZN(n480) );
  XNOR2_X1 U563 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U564 ( .A(n489), .B(n485), .ZN(n626) );
  NAND2_X1 U565 ( .A1(n626), .A2(n509), .ZN(n486) );
  XNOR2_X2 U566 ( .A(n486), .B(G472), .ZN(n682) );
  INV_X1 U567 ( .A(KEYINPUT105), .ZN(n487) );
  XNOR2_X1 U568 ( .A(n487), .B(KEYINPUT6), .ZN(n488) );
  XNOR2_X1 U569 ( .A(n682), .B(n488), .ZN(n590) );
  XNOR2_X1 U570 ( .A(KEYINPUT71), .B(G137), .ZN(n503) );
  NAND2_X1 U571 ( .A1(n731), .A2(G227), .ZN(n490) );
  XNOR2_X1 U572 ( .A(n490), .B(G140), .ZN(n492) );
  XNOR2_X1 U573 ( .A(KEYINPUT81), .B(G146), .ZN(n491) );
  XNOR2_X1 U574 ( .A(n492), .B(n491), .ZN(n493) );
  INV_X1 U575 ( .A(G469), .ZN(n495) );
  XNOR2_X2 U576 ( .A(n496), .B(n495), .ZN(n568) );
  XNOR2_X1 U577 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n497) );
  XNOR2_X2 U578 ( .A(n568), .B(n497), .ZN(n523) );
  NAND2_X1 U579 ( .A1(G221), .A2(n498), .ZN(n500) );
  XOR2_X1 U580 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n499) );
  XNOR2_X1 U581 ( .A(n500), .B(n499), .ZN(n507) );
  XOR2_X1 U582 ( .A(KEYINPUT87), .B(G110), .Z(n502) );
  XNOR2_X1 U583 ( .A(n502), .B(n501), .ZN(n505) );
  XNOR2_X1 U584 ( .A(n503), .B(KEYINPUT97), .ZN(n504) );
  XNOR2_X1 U585 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U586 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U587 ( .A(n508), .B(n729), .ZN(n632) );
  NAND2_X1 U588 ( .A1(n510), .A2(G217), .ZN(n512) );
  XNOR2_X1 U589 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n511) );
  XNOR2_X1 U590 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U591 ( .A1(n371), .A2(n674), .ZN(n514) );
  XOR2_X1 U592 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n515) );
  BUF_X1 U593 ( .A(n517), .Z(n518) );
  INV_X1 U594 ( .A(n518), .ZN(n521) );
  INV_X1 U595 ( .A(n674), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n682), .A2(n542), .ZN(n519) );
  NAND2_X1 U597 ( .A1(n523), .A2(n519), .ZN(n520) );
  NOR2_X1 U598 ( .A1(n521), .A2(n520), .ZN(n617) );
  OR2_X1 U599 ( .A1(n522), .A2(n674), .ZN(n677) );
  INV_X1 U600 ( .A(n590), .ZN(n524) );
  NAND2_X1 U601 ( .A1(n534), .A2(n699), .ZN(n525) );
  XNOR2_X1 U602 ( .A(n525), .B(KEYINPUT34), .ZN(n526) );
  NAND2_X1 U603 ( .A1(n538), .A2(n539), .ZN(n573) );
  NOR2_X2 U604 ( .A1(n526), .A2(n573), .ZN(n528) );
  XNOR2_X1 U605 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n527) );
  XNOR2_X2 U606 ( .A(n528), .B(n527), .ZN(n616) );
  NAND2_X1 U607 ( .A1(n546), .A2(n616), .ZN(n529) );
  INV_X1 U608 ( .A(n682), .ZN(n566) );
  NOR2_X1 U609 ( .A1(n530), .A2(n566), .ZN(n684) );
  NAND2_X1 U610 ( .A1(n534), .A2(n684), .ZN(n531) );
  XNOR2_X1 U611 ( .A(n531), .B(KEYINPUT31), .ZN(n665) );
  NOR2_X1 U612 ( .A1(n677), .A2(n568), .ZN(n533) );
  XNOR2_X1 U613 ( .A(n533), .B(n532), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n535), .A2(n682), .ZN(n652) );
  INV_X1 U615 ( .A(n539), .ZN(n536) );
  NOR2_X1 U616 ( .A1(n538), .A2(n536), .ZN(n537) );
  XNOR2_X1 U617 ( .A(KEYINPUT104), .B(n537), .ZN(n666) );
  INV_X1 U618 ( .A(n538), .ZN(n540) );
  XNOR2_X1 U619 ( .A(n541), .B(KEYINPUT90), .ZN(n543) );
  INV_X1 U620 ( .A(n616), .ZN(n544) );
  XNOR2_X1 U621 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n547) );
  XOR2_X1 U622 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n560) );
  NOR2_X1 U623 ( .A1(G900), .A2(n548), .ZN(n549) );
  NAND2_X1 U624 ( .A1(G953), .A2(n549), .ZN(n550) );
  XNOR2_X1 U625 ( .A(KEYINPUT107), .B(n550), .ZN(n551) );
  NOR2_X1 U626 ( .A1(n552), .A2(n551), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n682), .A2(n690), .ZN(n553) );
  XOR2_X1 U628 ( .A(KEYINPUT30), .B(n553), .Z(n554) );
  NAND2_X1 U629 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U630 ( .A1(n563), .A2(n556), .ZN(n575) );
  XOR2_X1 U631 ( .A(n600), .B(KEYINPUT38), .Z(n689) );
  NAND2_X1 U632 ( .A1(n575), .A2(n689), .ZN(n558) );
  XNOR2_X1 U633 ( .A(n558), .B(KEYINPUT39), .ZN(n596) );
  NAND2_X1 U634 ( .A1(n596), .A2(n663), .ZN(n559) );
  XNOR2_X1 U635 ( .A(n560), .B(n559), .ZN(n739) );
  INV_X1 U636 ( .A(n561), .ZN(n693) );
  NAND2_X1 U637 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U638 ( .A1(n693), .A2(n694), .ZN(n562) );
  XNOR2_X1 U639 ( .A(KEYINPUT41), .B(n562), .ZN(n707) );
  NOR2_X1 U640 ( .A1(n673), .A2(n563), .ZN(n564) );
  XOR2_X1 U641 ( .A(n564), .B(KEYINPUT73), .Z(n565) );
  XNOR2_X1 U642 ( .A(KEYINPUT28), .B(n567), .ZN(n570) );
  INV_X1 U643 ( .A(n568), .ZN(n569) );
  XNOR2_X1 U644 ( .A(n352), .B(KEYINPUT42), .ZN(n740) );
  NOR2_X1 U645 ( .A1(n739), .A2(n740), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n695), .A2(KEYINPUT47), .ZN(n572) );
  XNOR2_X1 U647 ( .A(n572), .B(KEYINPUT86), .ZN(n577) );
  INV_X1 U648 ( .A(n573), .ZN(n574) );
  AND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n576), .A2(n600), .ZN(n660) );
  NAND2_X1 U651 ( .A1(n577), .A2(n660), .ZN(n578) );
  XNOR2_X1 U652 ( .A(KEYINPUT85), .B(n578), .ZN(n585) );
  BUF_X1 U653 ( .A(n579), .Z(n580) );
  NAND2_X1 U654 ( .A1(KEYINPUT70), .A2(n661), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n581), .B(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n695), .A2(n661), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n594) );
  XOR2_X1 U659 ( .A(KEYINPUT92), .B(KEYINPUT36), .Z(n592) );
  INV_X1 U660 ( .A(n587), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n588), .A2(n663), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n586), .A2(n597), .ZN(n591) );
  XOR2_X1 U664 ( .A(n592), .B(n591), .Z(n593) );
  NOR2_X1 U665 ( .A1(n593), .A2(n523), .ZN(n668) );
  NOR2_X1 U666 ( .A1(n594), .A2(n668), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n666), .ZN(n670) );
  INV_X1 U668 ( .A(n670), .ZN(n603) );
  AND2_X1 U669 ( .A1(n597), .A2(n690), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n598), .A2(n523), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT43), .ZN(n602) );
  INV_X1 U672 ( .A(n600), .ZN(n601) );
  AND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n671) );
  NOR2_X1 U674 ( .A1(n603), .A2(n671), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT94), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT55), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n607), .B(n609), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U679 ( .A(G952), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n612), .A2(G953), .ZN(n635) );
  NAND2_X1 U681 ( .A1(n613), .A2(n635), .ZN(n615) );
  INV_X1 U682 ( .A(KEYINPUT56), .ZN(n614) );
  XNOR2_X1 U683 ( .A(n615), .B(n614), .ZN(G51) );
  XNOR2_X1 U684 ( .A(n616), .B(G122), .ZN(G24) );
  XOR2_X1 U685 ( .A(G110), .B(n617), .Z(G12) );
  XNOR2_X1 U686 ( .A(n618), .B(KEYINPUT59), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n621), .A2(n635), .ZN(n623) );
  XNOR2_X1 U689 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n622) );
  XNOR2_X1 U690 ( .A(n623), .B(n622), .ZN(G60) );
  XNOR2_X1 U691 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n624) );
  XOR2_X1 U692 ( .A(n624), .B(KEYINPUT62), .Z(n625) );
  XNOR2_X1 U693 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U694 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U695 ( .A1(n629), .A2(n635), .ZN(n630) );
  XNOR2_X1 U696 ( .A(n630), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U697 ( .A(n344), .B(G119), .Z(G21) );
  NAND2_X1 U698 ( .A1(n642), .A2(G217), .ZN(n634) );
  XNOR2_X1 U699 ( .A(n632), .B(KEYINPUT123), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(n636) );
  INV_X1 U701 ( .A(n635), .ZN(n647) );
  NOR2_X1 U702 ( .A1(n636), .A2(n647), .ZN(G66) );
  NAND2_X1 U703 ( .A1(n642), .A2(G478), .ZN(n640) );
  XNOR2_X1 U704 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X1 U707 ( .A1(n641), .A2(n647), .ZN(G63) );
  NAND2_X1 U708 ( .A1(n642), .A2(G469), .ZN(n646) );
  XOR2_X1 U709 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n643) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n646), .B(n645), .ZN(n648) );
  NOR2_X1 U712 ( .A1(n648), .A2(n647), .ZN(G54) );
  XOR2_X1 U713 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n650) );
  NAND2_X1 U714 ( .A1(n652), .A2(n663), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U716 ( .A(G104), .B(n651), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n654) );
  NAND2_X1 U718 ( .A1(n652), .A2(n666), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n654), .B(n653), .ZN(n656) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT113), .Z(n655) );
  XNOR2_X1 U721 ( .A(n656), .B(n655), .ZN(G9) );
  XOR2_X1 U722 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n658) );
  NAND2_X1 U723 ( .A1(n661), .A2(n666), .ZN(n657) );
  XNOR2_X1 U724 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U725 ( .A(G128), .B(n659), .ZN(G30) );
  XNOR2_X1 U726 ( .A(G143), .B(n660), .ZN(G45) );
  NAND2_X1 U727 ( .A1(n661), .A2(n663), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(G146), .ZN(G48) );
  NAND2_X1 U729 ( .A1(n665), .A2(n663), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(G113), .ZN(G15) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n667), .B(G116), .ZN(G18) );
  XNOR2_X1 U733 ( .A(n668), .B(G125), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U735 ( .A(G134), .B(n670), .ZN(G36) );
  XOR2_X1 U736 ( .A(G140), .B(n671), .Z(G42) );
  XNOR2_X1 U737 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT117), .ZN(n687) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n675), .B(KEYINPUT115), .ZN(n676) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(n676), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n523), .A2(n677), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(KEYINPUT50), .ZN(n679) );
  XNOR2_X1 U744 ( .A(KEYINPUT116), .B(n679), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U748 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U749 ( .A1(n707), .A2(n688), .ZN(n703) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U751 ( .A(KEYINPUT119), .B(n691), .Z(n692) );
  NOR2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n696), .B(KEYINPUT120), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n701) );
  INV_X1 U756 ( .A(n699), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U760 ( .A1(n706), .A2(n705), .ZN(n711) );
  INV_X1 U761 ( .A(n707), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n708), .A2(n699), .ZN(n709) );
  NAND2_X1 U763 ( .A1(n709), .A2(n731), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U767 ( .A(n715), .B(n716), .Z(n717) );
  XNOR2_X1 U768 ( .A(KEYINPUT125), .B(n717), .ZN(n719) );
  NOR2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n727) );
  OR2_X1 U770 ( .A1(n720), .A2(G953), .ZN(n725) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n722), .A2(G898), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(KEYINPUT126), .B(n728), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n730), .B(n733), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(n738) );
  XNOR2_X1 U780 ( .A(n733), .B(G227), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(G900), .ZN(n735) );
  XOR2_X1 U782 ( .A(KEYINPUT127), .B(n735), .Z(n736) );
  NAND2_X1 U783 ( .A1(G953), .A2(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U785 ( .A(G131), .B(n739), .Z(G33) );
  XOR2_X1 U786 ( .A(G137), .B(n740), .Z(G39) );
  XNOR2_X1 U787 ( .A(G101), .B(n741), .ZN(G3) );
endmodule

