//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n457), .B2(new_n458), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n473), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n473), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G124), .B2(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n476), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT70), .B1(new_n473), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n493), .A3(G2104), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n486), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n499), .A2(KEYINPUT72), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n500), .A2(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  XOR2_X1   g091(.A(KEYINPUT73), .B(G51), .Z(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(G89), .ZN(new_n520));
  OAI221_X1 g095(.A(new_n518), .B1(KEYINPUT7), .B2(new_n519), .C1(new_n513), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n506), .A2(G63), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n508), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G168));
  AOI22_X1  g100(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n508), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n511), .A2(G52), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n527), .A2(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  AOI22_X1  g107(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n508), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n511), .A2(G43), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n513), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT75), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G188));
  XNOR2_X1  g120(.A(KEYINPUT78), .B(G65), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n506), .A2(new_n546), .B1(G78), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n508), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n500), .A2(new_n502), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n504), .A2(new_n505), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n549), .A2(new_n550), .A3(new_n510), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G91), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n554));
  NAND3_X1  g129(.A1(new_n511), .A2(G53), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT77), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n511), .A2(new_n557), .A3(G53), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n511), .A2(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n551), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n511), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND4_X1  g144(.A1(new_n549), .A2(new_n550), .A3(G86), .A4(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n511), .A2(G48), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n549), .A2(new_n550), .A3(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT79), .B1(new_n576), .B2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n578));
  AOI211_X1 g153(.A(new_n578), .B(new_n508), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n572), .B(new_n573), .C1(new_n577), .C2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n508), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n511), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n513), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n551), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n589), .B(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n506), .A2(G66), .ZN(new_n596));
  INV_X1    g171(.A(G79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n501), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n592), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n562), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT82), .Z(G297));
  XOR2_X1   g180(.A(new_n604), .B(KEYINPUT83), .Z(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  INV_X1    g183(.A(new_n538), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n592), .A2(new_n595), .A3(new_n599), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(KEYINPUT84), .A3(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT84), .B1(new_n612), .B2(G559), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n611), .B1(new_n616), .B2(new_n610), .ZN(G323));
  XOR2_X1   g192(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n618));
  XNOR2_X1  g193(.A(G323), .B(new_n618), .ZN(G282));
  INV_X1    g194(.A(new_n477), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n620), .A2(KEYINPUT86), .A3(G135), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n477), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n482), .A2(G123), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n625), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n624), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT88), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n655), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n653), .A2(KEYINPUT17), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n662));
  OAI221_X1 g237(.A(new_n661), .B1(new_n659), .B2(new_n655), .C1(new_n662), .C2(new_n653), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n633), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2100), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(G2100), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  AOI22_X1  g253(.A1(new_n676), .A2(new_n677), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(new_n677), .C2(new_n676), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G29), .A2(G35), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G162), .B2(G29), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT29), .ZN(new_n691));
  INV_X1    g266(.A(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G26), .ZN(new_n695));
  OR3_X1    g270(.A1(KEYINPUT97), .A2(G104), .A3(G2105), .ZN(new_n696));
  INV_X1    g271(.A(G116), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n462), .B1(new_n697), .B2(G2105), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT97), .B1(G104), .B2(G2105), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT98), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n482), .A2(G128), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n620), .A2(G140), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT99), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n695), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  MUX2_X1   g283(.A(new_n695), .B(new_n708), .S(KEYINPUT28), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT100), .B(G2067), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G28), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(G28), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n713), .A2(new_n714), .A3(G29), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT101), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G33), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n716), .A2(G29), .A3(G33), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n620), .A2(G139), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n721), .C1(new_n473), .C2(new_n722), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n717), .B(new_n718), .C1(new_n723), .C2(new_n694), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G2072), .Z(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G32), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n476), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G2105), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n728), .B(new_n730), .C1(G129), .C2(new_n482), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT27), .B(G1996), .Z(new_n733));
  AOI211_X1 g308(.A(new_n715), .B(new_n725), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n735), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1966), .ZN(new_n738));
  NOR2_X1   g313(.A1(G27), .A2(G29), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G164), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT103), .B(G2078), .Z(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G11), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n632), .A2(new_n694), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n734), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n735), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n735), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1961), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n740), .B2(new_n741), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(G1961), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT95), .B(G16), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT104), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1956), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n694), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n694), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n753), .A2(G19), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n538), .B2(new_n753), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G1341), .Z(new_n768));
  NAND4_X1  g343(.A1(new_n751), .A2(new_n758), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n711), .A2(new_n745), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n694), .A2(G25), .ZN(new_n771));
  INV_X1    g346(.A(G131), .ZN(new_n772));
  OR3_X1    g347(.A1(new_n477), .A2(KEYINPUT92), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n477), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n482), .A2(G119), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT93), .Z(new_n779));
  AOI21_X1  g354(.A(new_n771), .B1(new_n779), .B2(G29), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n771), .B(new_n780), .S(KEYINPUT91), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT35), .B(G1991), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT94), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n752), .A2(G24), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n586), .B2(new_n752), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G1986), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G1986), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n753), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n753), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT96), .Z(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1971), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G1971), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1976), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n735), .A2(G6), .ZN(new_n801));
  INV_X1    g376(.A(G305), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n735), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n795), .A2(KEYINPUT34), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n800), .A2(new_n793), .A3(new_n794), .ZN(new_n808));
  INV_X1    g383(.A(new_n805), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n789), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n789), .B2(new_n811), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n693), .B(new_n770), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n735), .A2(G4), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n600), .B2(new_n735), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1348), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n732), .A2(new_n733), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT102), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n815), .A2(new_n818), .A3(new_n820), .ZN(G311));
  INV_X1    g396(.A(new_n770), .ZN(new_n822));
  INV_X1    g397(.A(new_n814), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n789), .A2(new_n811), .A3(new_n812), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n818), .ZN(new_n826));
  INV_X1    g401(.A(new_n820), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n693), .ZN(G150));
  AOI22_X1  g403(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n508), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n511), .A2(G55), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n513), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n538), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n612), .A2(new_n607), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n844), .B2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT105), .ZN(G145));
  XNOR2_X1  g421(.A(new_n779), .B(KEYINPUT107), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n706), .B(new_n622), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n731), .B(new_n723), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n632), .B(G160), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G162), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n482), .A2(G130), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n620), .A2(G142), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n496), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n853), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n851), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n851), .A2(new_n862), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g442(.A1(new_n615), .A2(new_n840), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n838), .A2(new_n839), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n613), .B2(new_n614), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n600), .A2(new_n562), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n612), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(KEYINPUT41), .A3(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OAI22_X1  g453(.A1(new_n868), .A2(new_n870), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n871), .A2(new_n872), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n868), .A2(new_n881), .A3(new_n870), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G166), .B(G288), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G305), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  INV_X1    g463(.A(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n879), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n883), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n883), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(G868), .B2(new_n834), .ZN(G331));
  XNOR2_X1  g471(.A(new_n840), .B(G286), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G171), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n869), .A2(G286), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n840), .A2(G168), .ZN(new_n900));
  OAI21_X1  g475(.A(G301), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n876), .B2(new_n878), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n873), .A3(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n886), .A3(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n898), .A2(new_n901), .B1(new_n875), .B2(new_n877), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n898), .A2(new_n873), .A3(new_n901), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n887), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n908), .A3(new_n864), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n905), .A2(new_n908), .A3(new_n911), .A4(new_n864), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(G397));
  NOR2_X1   g490(.A1(new_n706), .A2(G2067), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n706), .A2(G2067), .ZN(new_n918));
  INV_X1    g493(.A(G1996), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n731), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n496), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n469), .A2(new_n474), .A3(G40), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n919), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT109), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n920), .A2(new_n926), .B1(new_n731), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n779), .A2(new_n783), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n779), .A2(new_n783), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n586), .B(G1986), .Z(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT122), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT49), .ZN(new_n937));
  INV_X1    g512(.A(G1981), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n578), .B1(new_n939), .B2(new_n508), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n576), .A2(KEYINPUT79), .A3(G651), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n940), .A2(new_n941), .B1(G48), .B2(new_n511), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n942), .B2(new_n570), .ZN(new_n943));
  NOR2_X1   g518(.A1(G305), .A2(G1981), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G8), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n469), .A2(new_n474), .A3(G40), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n496), .A2(new_n921), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n573), .B1(new_n577), .B2(new_n579), .ZN(new_n950));
  INV_X1    g525(.A(new_n570), .ZN(new_n951));
  OAI21_X1  g526(.A(G1981), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n945), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n496), .B2(new_n921), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n956), .A2(new_n957), .A3(new_n925), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n958), .B2(G1971), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n922), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n496), .A2(KEYINPUT50), .A3(new_n921), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n925), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n692), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n924), .A2(new_n947), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1971), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n509), .B2(new_n515), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(G8), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n970), .B(KEYINPUT55), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n692), .A2(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n946), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(G1976), .ZN(new_n977));
  AND2_X1   g552(.A1(G288), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(new_n978), .B2(new_n949), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n566), .A2(G1976), .A3(new_n567), .A4(new_n568), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n949), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n981), .B(new_n949), .C1(new_n978), .C2(KEYINPUT52), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n954), .A2(new_n973), .A3(new_n976), .A4(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n496), .A2(KEYINPUT50), .A3(new_n921), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT50), .B1(new_n496), .B2(new_n921), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n947), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1961), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT117), .B(new_n947), .C1(new_n987), .C2(new_n988), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n966), .A2(new_n995), .A3(G2078), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n966), .B2(G2078), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n996), .A3(G301), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(KEYINPUT54), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n986), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n989), .B2(G2084), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n966), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n961), .A2(new_n962), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT113), .A3(new_n764), .A4(new_n947), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G286), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1008), .A2(new_n1013), .A3(new_n1009), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(G8), .C1(new_n1007), .C2(G286), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(G8), .A3(G286), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT54), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(G171), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(G171), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(new_n1020), .A3(KEYINPUT54), .A4(new_n998), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1000), .A2(new_n1018), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(G1348), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n991), .A2(new_n1027), .A3(new_n993), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n947), .A2(new_n948), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(G2067), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1026), .B1(new_n1033), .B2(new_n600), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT60), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(KEYINPUT119), .A3(new_n612), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1034), .A2(new_n1036), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n553), .B2(new_n561), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n556), .A2(new_n560), .A3(new_n558), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(new_n548), .A3(KEYINPUT57), .A4(new_n552), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n958), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1956), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n989), .A2(KEYINPUT115), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT115), .B1(new_n989), .B2(new_n1045), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1042), .B(new_n1044), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1048), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1046), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT116), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT58), .B(G1341), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1029), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(G1996), .B2(new_n966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n538), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT59), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1063), .B(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1049), .A2(KEYINPUT61), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(new_n1053), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1033), .A2(new_n1026), .A3(new_n600), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n1035), .B2(new_n612), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1037), .A2(new_n1059), .A3(new_n1069), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1042), .B1(new_n1055), .B2(new_n1044), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n600), .B2(new_n1031), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1025), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n969), .A2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n974), .A2(KEYINPUT114), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1007), .A2(G8), .A3(G168), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n954), .B(new_n985), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT63), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n954), .A2(new_n1089), .A3(new_n797), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n949), .B1(new_n1090), .B2(new_n944), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n976), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n973), .B1(new_n1093), .B2(new_n1084), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n954), .A3(new_n985), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n936), .B1(new_n1080), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1096), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1071), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1063), .B1(new_n1064), .B2(KEYINPUT59), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1065), .B1(new_n1062), .B2(new_n538), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1067), .A2(new_n1075), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1078), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT122), .B(new_n1098), .C1(new_n1106), .C2(new_n1025), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1018), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n986), .A2(new_n1023), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1014), .A2(new_n1016), .A3(new_n1115), .A4(new_n1017), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1114), .A2(KEYINPUT123), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT123), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT125), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1113), .B(new_n1121), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n935), .B1(new_n1108), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n928), .B(KEYINPUT46), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n917), .A2(new_n731), .A3(new_n918), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n926), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n916), .B1(new_n929), .B2(new_n931), .ZN(new_n1129));
  INV_X1    g704(.A(new_n926), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(G1986), .A3(G290), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT126), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT48), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1129), .A2(new_n1130), .B1(new_n933), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g711(.A1(new_n666), .A2(G319), .A3(new_n667), .ZN(new_n1138));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n1139));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1141));
  NOR3_X1   g715(.A1(G401), .A2(G229), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g716(.A1(new_n913), .A2(new_n866), .A3(new_n1140), .A4(new_n1142), .ZN(G225));
  INV_X1    g717(.A(G225), .ZN(G308));
endmodule


