//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879;
  XNOR2_X1  g000(.A(KEYINPUT85), .B(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n209), .C1(KEYINPUT15), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G1gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT88), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n218), .B(new_n219), .C1(G1gat), .C2(new_n216), .ZN(new_n220));
  INV_X1    g019(.A(G8gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n213), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT89), .B1(new_n224), .B2(new_n225), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(new_n226), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n228), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n228), .A3(new_n226), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G141gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT83), .ZN(new_n239));
  XOR2_X1   g038(.A(G169gat), .B(G197gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n229), .A2(new_n245), .A3(new_n233), .A4(new_n236), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(KEYINPUT90), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G120gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT1), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G127gat), .B(G134gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT70), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT1), .B1(new_n264), .B2(KEYINPUT69), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n257), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n259), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G141gat), .B(G148gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT2), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n276), .B(new_n275), .C1(new_n271), .C2(KEYINPUT2), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n270), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n270), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n269), .B1(new_n261), .B2(new_n262), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n281), .ZN(new_n292));
  AND2_X1   g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n284), .A2(new_n290), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n282), .A2(new_n293), .ZN(new_n296));
  AND4_X1   g095(.A1(new_n284), .A2(new_n296), .A3(new_n290), .A4(new_n292), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n263), .A2(new_n270), .A3(new_n281), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n281), .B1(new_n263), .B2(new_n270), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT0), .B(G57gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(G85gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n295), .C1(new_n297), .C2(new_n301), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n302), .A2(KEYINPUT6), .A3(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G64gat), .ZN(new_n315));
  INV_X1    g114(.A(G92gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT26), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(KEYINPUT26), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n323), .B(new_n324), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(KEYINPUT28), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT28), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n329), .B(new_n330), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  AND2_X1   g137(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n340));
  OAI211_X1 g139(.A(KEYINPUT23), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT24), .A3(new_n330), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n330), .A2(KEYINPUT24), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n326), .A2(new_n328), .B1(KEYINPUT23), .B2(new_n321), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n337), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n325), .A2(G169gat), .A3(G176gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n349), .A2(new_n322), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n321), .B2(KEYINPUT23), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n352), .A2(new_n343), .A3(new_n344), .A4(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n347), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n347), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n336), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT74), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n336), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n320), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT72), .B(G218gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT22), .B1(new_n363), .B2(G211gat), .ZN(new_n364));
  XOR2_X1   g163(.A(G197gat), .B(G204gat), .Z(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n366), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n355), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n336), .A2(new_n370), .A3(new_n318), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n362), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n318), .A3(new_n361), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n336), .A2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n319), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n379), .A2(KEYINPUT37), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(KEYINPUT37), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n317), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n313), .B1(new_n382), .B2(KEYINPUT38), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n377), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n369), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n347), .A2(new_n348), .A3(new_n355), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n360), .B1(new_n388), .B2(new_n336), .ZN(new_n389));
  INV_X1    g188(.A(new_n361), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n319), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n374), .A3(new_n371), .ZN(new_n392));
  INV_X1    g191(.A(new_n317), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT38), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n369), .B1(new_n362), .B2(new_n372), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n374), .A3(new_n377), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(KEYINPUT37), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(new_n317), .C1(new_n381), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n366), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n403), .B(new_n404), .C1(new_n366), .C2(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n281), .B1(new_n405), .B2(new_n288), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n369), .B1(new_n404), .B2(new_n289), .ZN(new_n407));
  INV_X1    g206(.A(G228gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  OAI22_X1  g208(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n289), .A2(new_n404), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n374), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n408), .A2(new_n409), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n369), .B2(new_n404), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n281), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G22gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G78gat), .ZN(new_n424));
  INV_X1    g223(.A(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n421), .A2(new_n418), .A3(new_n417), .A4(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n421), .A2(new_n417), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n419), .B(new_n427), .C1(new_n428), .C2(new_n426), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n284), .A2(new_n290), .A3(new_n292), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n293), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n298), .A2(new_n299), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(KEYINPUT39), .C1(new_n293), .C2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n306), .C1(KEYINPUT39), .C2(new_n432), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n437), .B(KEYINPUT40), .Z(new_n438));
  NAND4_X1  g237(.A1(new_n379), .A2(KEYINPUT75), .A3(KEYINPUT30), .A4(new_n393), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n385), .A2(new_n392), .A3(KEYINPUT30), .A4(new_n393), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n393), .B1(new_n385), .B2(new_n392), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n394), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n447), .A3(new_n308), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n400), .A2(new_n430), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n358), .A2(new_n285), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n291), .B(new_n336), .C1(new_n356), .C2(new_n357), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G227gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n409), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT64), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n450), .B(new_n451), .C1(new_n454), .C2(new_n409), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G15gat), .B(G43gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n456), .B1(new_n450), .B2(new_n451), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(KEYINPUT33), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI221_X4 g269(.A(new_n468), .B1(KEYINPUT33), .B2(new_n465), .C1(new_n452), .C2(new_n457), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n291), .B1(new_n388), .B2(new_n336), .ZN(new_n473));
  INV_X1    g272(.A(new_n451), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n478), .A3(new_n465), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n467), .A2(new_n469), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n453), .A2(new_n458), .B1(new_n460), .B2(KEYINPUT34), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n472), .A2(KEYINPUT71), .A3(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n462), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n311), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n309), .A4(new_n310), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n312), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n443), .A2(new_n495), .A3(new_n446), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n449), .B(new_n491), .C1(new_n496), .C2(new_n430), .ZN(new_n497));
  INV_X1    g296(.A(new_n447), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n429), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n313), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n429), .B1(new_n486), .B2(new_n488), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT81), .B1(new_n503), .B2(KEYINPUT35), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n505), .B(new_n499), .C1(new_n496), .C2(new_n502), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n253), .B1(new_n497), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509));
  INV_X1    g308(.A(G71gat), .ZN(new_n510));
  INV_X1    g309(.A(G78gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT92), .ZN(new_n515));
  XOR2_X1   g314(.A(G57gat), .B(G64gat), .Z(new_n516));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n517), .A3(new_n513), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n516), .A2(KEYINPUT9), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT91), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n513), .A3(new_n524), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n222), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G183gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G127gat), .B(G155gat), .ZN(new_n533));
  INV_X1    g332(.A(G211gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n526), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n537), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n532), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G190gat), .B(G218gat), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT100), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n544), .B1(new_n545), .B2(new_n316), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT98), .Z(new_n554));
  AND2_X1   g353(.A1(new_n215), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n213), .B2(new_n553), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT99), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n543), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n542), .A2(KEYINPUT100), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT96), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n560), .B(new_n562), .Z(new_n563));
  AND2_X1   g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n559), .A2(new_n563), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n553), .B(new_n526), .Z(new_n570));
  INV_X1    g369(.A(KEYINPUT10), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n553), .A2(new_n526), .A3(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n570), .A2(new_n575), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G120gat), .B(G148gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G176gat), .ZN(new_n580));
  INV_X1    g379(.A(G204gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  AND4_X1   g382(.A1(new_n541), .A2(new_n568), .A3(new_n569), .A4(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n508), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n495), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT101), .B(G1gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(G1324gat));
  AND2_X1   g388(.A1(new_n585), .A2(new_n447), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n217), .A2(new_n221), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT42), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(KEYINPUT42), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n594), .B(new_n595), .C1(new_n221), .C2(new_n590), .ZN(G1325gat));
  AOI21_X1  g395(.A(G15gat), .B1(new_n585), .B2(new_n484), .ZN(new_n597));
  INV_X1    g396(.A(new_n491), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(G15gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n585), .B2(new_n599), .ZN(G1326gat));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n429), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT43), .B(G22gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(G1327gat));
  NAND2_X1  g402(.A1(new_n568), .A2(new_n569), .ZN(new_n604));
  INV_X1    g403(.A(new_n583), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n541), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n508), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n607), .A2(new_n495), .A3(new_n202), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT45), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n507), .A2(KEYINPUT102), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n611), .B(new_n501), .C1(new_n504), .C2(new_n506), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n497), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n604), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n604), .ZN(new_n617));
  AOI211_X1 g416(.A(new_n615), .B(new_n617), .C1(new_n497), .C2(new_n507), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n616), .A2(new_n249), .A3(new_n606), .A4(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n202), .B1(new_n620), .B2(new_n495), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n609), .A2(new_n621), .ZN(G1328gat));
  OR2_X1    g421(.A1(new_n498), .A2(G36gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT46), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(KEYINPUT46), .ZN(new_n629));
  OAI21_X1  g428(.A(G36gat), .B1(new_n620), .B2(new_n498), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n626), .B2(KEYINPUT46), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(G1329gat));
  INV_X1    g431(.A(G43gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n607), .B2(new_n483), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n491), .A2(new_n633), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n634), .B(new_n635), .C1(new_n620), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT106), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n618), .B1(new_n614), .B2(new_n615), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n640), .A2(new_n249), .A3(new_n606), .A4(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT47), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n641), .A2(new_n644), .A3(new_n634), .A4(new_n635), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n639), .A2(new_n643), .A3(new_n648), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(G1330gat));
  NAND2_X1  g449(.A1(new_n429), .A2(G50gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n607), .A2(new_n430), .ZN(new_n652));
  OAI22_X1  g451(.A1(new_n620), .A2(new_n651), .B1(G50gat), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g453(.A(new_n249), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n613), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n541), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n656), .A2(new_n657), .A3(new_n604), .A4(new_n583), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n586), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g459(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n447), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(KEYINPUT108), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(KEYINPUT108), .ZN(new_n664));
  OR2_X1    g463(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n663), .B2(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1333gat));
  AOI21_X1  g467(.A(new_n510), .B1(new_n658), .B2(new_n598), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n658), .A2(new_n510), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n484), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g471(.A1(new_n658), .A2(new_n429), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT109), .B(G78gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1335gat));
  NOR2_X1   g474(.A1(new_n249), .A2(new_n541), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n605), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n640), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G85gat), .B1(new_n679), .B2(new_n495), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n613), .A2(new_n604), .A3(new_n676), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT51), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n605), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n586), .A2(new_n545), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT110), .ZN(G1336gat));
  NAND3_X1  g486(.A1(new_n447), .A2(new_n605), .A3(new_n316), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT111), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT52), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n640), .A2(new_n447), .A3(new_n678), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT113), .ZN(new_n693));
  OAI21_X1  g492(.A(G92gat), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n677), .B(new_n618), .C1(new_n614), .C2(new_n615), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT113), .B1(new_n695), .B2(new_n447), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n691), .B(KEYINPUT114), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(KEYINPUT113), .A3(new_n447), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(G92gat), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT114), .B1(new_n701), .B2(new_n691), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n682), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT112), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n681), .B(KEYINPUT51), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(KEYINPUT112), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(new_n690), .B1(G92gat), .B2(new_n692), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n698), .A2(new_n702), .B1(new_n703), .B2(new_n708), .ZN(G1337gat));
  OAI21_X1  g508(.A(G99gat), .B1(new_n679), .B2(new_n491), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n483), .A2(G99gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n684), .B2(new_n711), .ZN(G1338gat));
  OAI21_X1  g511(.A(G106gat), .B1(new_n679), .B2(new_n430), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n605), .A2(new_n425), .A3(new_n429), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n713), .B(new_n714), .C1(new_n706), .C2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(KEYINPUT115), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(new_n713), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(new_n714), .ZN(G1339gat));
  INV_X1    g519(.A(new_n582), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT54), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n576), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT54), .B1(new_n574), .B2(new_n575), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n723), .B(KEYINPUT55), .C1(new_n576), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n578), .A2(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n576), .B2(new_n724), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n249), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n227), .A2(new_n228), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n231), .A2(new_n232), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n243), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n248), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(new_n605), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n617), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n604), .A2(new_n735), .A3(new_n730), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n541), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n584), .A2(new_n655), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n495), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n502), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n447), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n256), .A3(new_n249), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n739), .A2(new_n740), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n447), .A2(new_n495), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n500), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G113gat), .B1(new_n748), .B2(new_n253), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(G1340gat));
  NAND3_X1  g549(.A1(new_n744), .A2(new_n254), .A3(new_n605), .ZN(new_n751));
  OAI21_X1  g550(.A(G120gat), .B1(new_n748), .B2(new_n583), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1341gat));
  INV_X1    g552(.A(G127gat), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n748), .A2(new_n754), .A3(new_n657), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n541), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n754), .ZN(G1342gat));
  NOR2_X1   g556(.A1(new_n743), .A2(G134gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n604), .A2(new_n498), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT116), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT56), .Z(new_n762));
  OAI21_X1  g561(.A(G134gat), .B1(new_n748), .B2(new_n617), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1343gat));
  NAND3_X1  g563(.A1(new_n491), .A2(KEYINPUT120), .A3(new_n429), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n598), .B2(new_n430), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n253), .A2(G141gat), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(KEYINPUT121), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(KEYINPUT121), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n768), .A2(new_n447), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(KEYINPUT58), .ZN(new_n773));
  INV_X1    g572(.A(new_n727), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n729), .A2(KEYINPUT118), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT118), .B1(new_n729), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n774), .B(KEYINPUT119), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n251), .A2(new_n252), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n736), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n604), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n738), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n657), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n429), .B1(new_n787), .B2(new_n740), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT57), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n491), .A2(new_n747), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n741), .A2(new_n430), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G141gat), .B1(new_n794), .B2(new_n253), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n773), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n789), .A2(new_n249), .A3(new_n790), .A4(new_n793), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n772), .B1(new_n798), .B2(G141gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1344gat));
  NOR2_X1   g599(.A1(new_n768), .A2(new_n447), .ZN(new_n801));
  INV_X1    g600(.A(G148gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n605), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n804), .B(G148gat), .C1(new_n794), .C2(new_n583), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n792), .B1(new_n746), .B2(new_n429), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n584), .A2(new_n253), .A3(KEYINPUT122), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT122), .B1(new_n584), .B2(new_n253), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT57), .B(new_n430), .C1(new_n786), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n605), .A3(new_n790), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n804), .B1(new_n813), .B2(G148gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n803), .B1(new_n806), .B2(new_n814), .ZN(G1345gat));
  AOI21_X1  g614(.A(G155gat), .B1(new_n801), .B2(new_n541), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n794), .A2(new_n273), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n541), .ZN(G1346gat));
  OAI21_X1  g617(.A(G162gat), .B1(new_n794), .B2(new_n617), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n760), .A2(new_n274), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n768), .B2(new_n820), .ZN(G1347gat));
  NOR2_X1   g620(.A1(new_n498), .A2(new_n586), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n746), .A2(new_n502), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n338), .A3(new_n249), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT123), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n746), .A2(new_n500), .A3(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT124), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n746), .A2(new_n829), .A3(new_n500), .A4(new_n822), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G169gat), .B1(new_n831), .B2(new_n253), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(G1348gat));
  NOR4_X1   g632(.A1(new_n831), .A2(new_n340), .A3(new_n339), .A4(new_n583), .ZN(new_n834));
  AOI21_X1  g633(.A(G176gat), .B1(new_n824), .B2(new_n605), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1349gat));
  OAI21_X1  g635(.A(G183gat), .B1(new_n831), .B2(new_n657), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n824), .A2(new_n331), .A3(new_n541), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n828), .A2(new_n604), .A3(new_n830), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(G190gat), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n842), .B2(G190gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n842), .A2(G190gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT125), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(KEYINPUT61), .A3(new_n844), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n824), .A2(new_n332), .A3(new_n604), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(G1351gat));
  AND2_X1   g651(.A1(new_n491), .A2(new_n822), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n791), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n249), .ZN(new_n855));
  INV_X1    g654(.A(G197gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT126), .B1(new_n807), .B2(new_n811), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n786), .A2(new_n810), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n792), .A3(new_n429), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n860), .B(new_n861), .C1(new_n792), .C2(new_n791), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n858), .A2(new_n862), .A3(G197gat), .A4(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n857), .B1(new_n863), .B2(new_n253), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT127), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT127), .B(new_n857), .C1(new_n863), .C2(new_n253), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1352gat));
  NAND3_X1  g667(.A1(new_n854), .A2(new_n581), .A3(new_n605), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT62), .Z(new_n870));
  AND4_X1   g669(.A1(new_n605), .A2(new_n858), .A3(new_n862), .A4(new_n853), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n581), .B2(new_n871), .ZN(G1353gat));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n534), .A3(new_n541), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n812), .A2(new_n541), .A3(new_n853), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT63), .B1(new_n874), .B2(G211gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(G1354gat));
  AOI21_X1  g676(.A(G218gat), .B1(new_n854), .B2(new_n604), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n604), .A2(new_n858), .A3(new_n862), .A4(new_n853), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n363), .ZN(G1355gat));
endmodule


