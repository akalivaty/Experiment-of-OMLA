//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G224), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT87), .Z(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT7), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  AND4_X1   g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .A4(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n197), .A2(G128), .B1(new_n193), .B2(new_n195), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT0), .B(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n193), .A2(new_n195), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(KEYINPUT0), .A3(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n201), .A2(new_n202), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n190), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT2), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT2), .A2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G116), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n218), .A2(new_n222), .A3(new_n224), .A4(new_n219), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(KEYINPUT68), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT80), .A3(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(new_n232), .A3(KEYINPUT80), .A4(G104), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(G104), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(G101), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n234), .A2(new_n238), .A3(new_n243), .A4(new_n236), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n231), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT5), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(G113), .C1(KEYINPUT5), .C2(new_n222), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n227), .ZN(new_n249));
  INV_X1    g063(.A(G104), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G107), .ZN(new_n251));
  OAI21_X1  g065(.A(G101), .B1(new_n251), .B2(new_n237), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G122), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n246), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(KEYINPUT8), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n249), .A2(new_n253), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n214), .A2(KEYINPUT7), .A3(new_n189), .A4(new_n201), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n217), .A2(new_n257), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n255), .ZN(new_n265));
  INV_X1    g079(.A(new_n256), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n267), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n257), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n214), .A2(new_n201), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n269), .B(new_n189), .Z(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G210), .B1(G237), .B2(G902), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n264), .A2(new_n273), .A3(new_n275), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(KEYINPUT89), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n278), .A2(KEYINPUT89), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G214), .B1(G237), .B2(G902), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT85), .Z(new_n283));
  OAI21_X1  g097(.A(KEYINPUT90), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  INV_X1    g099(.A(new_n283), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n279), .A2(new_n280), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT9), .B(G234), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G221), .B1(new_n290), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G227), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G953), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n293), .B(new_n295), .Z(new_n296));
  INV_X1    g110(.A(KEYINPUT81), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n253), .B2(new_n199), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n197), .A2(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n208), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n205), .A2(G128), .A3(new_n197), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(KEYINPUT81), .A3(new_n244), .A4(new_n252), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT65), .A4(new_n312), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(G131), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n309), .A2(new_n311), .A3(new_n318), .A4(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n313), .B2(new_n314), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT66), .A3(new_n316), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n207), .A2(new_n211), .A3(new_n212), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n245), .A2(new_n326), .A3(new_n241), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n244), .A2(new_n252), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT10), .A3(new_n302), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n306), .A2(new_n325), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n329), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT10), .B1(new_n298), .B2(new_n303), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT82), .A3(new_n325), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n298), .A2(new_n303), .B1(new_n199), .B2(new_n253), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n325), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n338), .A2(new_n325), .A3(KEYINPUT12), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n296), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n335), .A2(new_n325), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT82), .B1(new_n335), .B2(new_n325), .ZN(new_n346));
  NOR4_X1   g160(.A1(new_n333), .A2(new_n334), .A3(new_n331), .A4(new_n324), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n296), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n345), .B1(new_n348), .B2(KEYINPUT83), .ZN(new_n349));
  INV_X1    g163(.A(new_n296), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n332), .B2(new_n336), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n344), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G469), .B1(new_n354), .B2(G902), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n337), .A2(new_n343), .A3(new_n296), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n351), .A2(KEYINPUT84), .A3(new_n343), .ZN(new_n359));
  INV_X1    g173(.A(new_n345), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n337), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n350), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G469), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT72), .B(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n292), .B1(new_n355), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n288), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n366), .B2(G234), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n221), .A2(G128), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n374));
  INV_X1    g188(.A(G128), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(G119), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n221), .A2(KEYINPUT23), .A3(G128), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT24), .B(G110), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n378), .A2(G110), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT74), .A2(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G140), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT74), .A3(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT16), .B1(new_n387), .B2(G125), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n192), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n386), .B2(new_n388), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n395), .A2(G146), .A3(new_n391), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n384), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(new_n192), .A3(new_n392), .ZN(new_n400));
  OAI21_X1  g214(.A(G146), .B1(new_n395), .B2(new_n391), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT75), .A3(new_n384), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n380), .A2(new_n382), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT76), .B(G110), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n373), .C1(new_n376), .C2(new_n377), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n380), .A2(new_n382), .A3(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n192), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n404), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n411), .A2(new_n414), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n399), .B2(new_n403), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT22), .B(G137), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n420), .B2(KEYINPUT79), .ZN(new_n427));
  AOI211_X1 g241(.A(new_n417), .B(new_n419), .C1(new_n399), .C2(new_n403), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT25), .B1(new_n430), .B2(new_n366), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n432), .B(new_n365), .C1(new_n426), .C2(new_n429), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n372), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n372), .A2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT28), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n213), .B1(new_n321), .B2(new_n323), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n319), .A2(KEYINPUT67), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n310), .A2(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n312), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(KEYINPUT67), .A3(G131), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n302), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n231), .B1(new_n440), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n322), .A2(KEYINPUT66), .A3(new_n316), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n322), .A2(new_n316), .B1(KEYINPUT66), .B2(new_n319), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n326), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n231), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n439), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n454), .A2(new_n439), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G237), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n187), .A3(G210), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n243), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n460), .B(new_n461), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT71), .B1(new_n457), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n365), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n440), .B2(new_n448), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n447), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n231), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n473), .A2(new_n454), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n464), .B1(new_n474), .B2(new_n462), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n453), .B1(new_n452), .B2(new_n447), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT69), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n439), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n449), .A2(new_n454), .A3(KEYINPUT69), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n456), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n475), .B1(new_n462), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G472), .B1(new_n469), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(new_n462), .A3(new_n454), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT31), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT31), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n473), .A2(new_n485), .A3(new_n462), .A4(new_n454), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n484), .B(new_n486), .C1(new_n462), .C2(new_n480), .ZN(new_n487));
  NOR2_X1   g301(.A1(G472), .A2(G902), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT73), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n484), .A2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n478), .A2(new_n479), .ZN(new_n492));
  INV_X1    g306(.A(new_n456), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n462), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n488), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(new_n497), .A3(new_n488), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT32), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT73), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n489), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n482), .B(new_n490), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n458), .A2(new_n187), .A3(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n194), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n458), .A2(new_n187), .A3(G143), .A4(G214), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n318), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(KEYINPUT18), .A3(G131), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n389), .A2(G146), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n413), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(G131), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT91), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n402), .B1(new_n517), .B2(KEYINPUT17), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n516), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n318), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n515), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n250), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n263), .B1(new_n524), .B2(new_n527), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n520), .A2(new_n522), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n535));
  AOI22_X1  g349(.A1(new_n412), .A2(new_n535), .B1(new_n389), .B2(KEYINPUT19), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n192), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n401), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n526), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n514), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n532), .A2(new_n533), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n540), .B(new_n541), .C1(new_n524), .C2(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT20), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n530), .A2(G475), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(G234), .A2(G237), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G952), .A3(new_n187), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n365), .A2(G953), .A3(new_n546), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT21), .B(G898), .Z(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n223), .A2(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n223), .A2(G122), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G107), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n232), .ZN(new_n556));
  XNOR2_X1  g370(.A(G128), .B(G143), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n308), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n559), .A2(new_n375), .A3(G143), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n560), .A2(KEYINPUT94), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(KEYINPUT94), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n194), .A2(G128), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT13), .B1(new_n194), .B2(G128), .ZN(new_n564));
  NOR4_X1   g378(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n558), .B1(new_n565), .B2(new_n308), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n556), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n557), .B(new_n308), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n553), .A2(KEYINPUT14), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n552), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n553), .A2(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g386(.A(G107), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n556), .A2(new_n567), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n569), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n290), .A2(new_n371), .A3(G953), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n566), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n566), .B2(new_n575), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n365), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT15), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n581), .A2(KEYINPUT96), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(KEYINPUT96), .ZN(new_n583));
  OAI21_X1  g397(.A(G478), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n580), .B(new_n584), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n551), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n370), .A2(new_n438), .A3(new_n503), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n487), .B2(new_n366), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n496), .B2(new_n498), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n368), .A2(new_n438), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n530), .A2(G475), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n542), .A2(new_n544), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n580), .A2(G478), .ZN(new_n597));
  AND2_X1   g411(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n598));
  NOR2_X1   g412(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n579), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n598), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n577), .B2(new_n578), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n600), .A2(G478), .A3(new_n366), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n283), .B1(new_n277), .B2(new_n278), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n550), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n593), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT34), .B(G104), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  OR2_X1    g425(.A1(new_n544), .A2(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT98), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n612), .A2(new_n594), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n614), .A2(new_n586), .A3(new_n550), .A4(new_n607), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n593), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT35), .B(G107), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  INV_X1    g432(.A(new_n372), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n427), .A2(new_n428), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n416), .A2(new_n417), .A3(new_n425), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n366), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n432), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n430), .A2(KEYINPUT25), .A3(new_n366), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n425), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n416), .B(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n435), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT99), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  INV_X1    g446(.A(new_n630), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n434), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n587), .A2(new_n592), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n369), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  INV_X1    g452(.A(new_n368), .ZN(new_n639));
  INV_X1    g453(.A(new_n607), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n631), .A2(new_n634), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  OR3_X1    g457(.A1(new_n548), .A2(new_n643), .A3(G900), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n548), .B2(G900), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n547), .B(KEYINPUT101), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT102), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n614), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n585), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n642), .A2(new_n503), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XOR2_X1   g468(.A(new_n649), .B(KEYINPUT39), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n368), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n641), .A2(new_n586), .A3(new_n596), .A4(new_n286), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n281), .B(KEYINPUT38), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n474), .A2(new_n463), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n449), .A2(new_n454), .A3(new_n463), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n263), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT103), .Z(new_n665));
  OAI211_X1 g479(.A(new_n490), .B(new_n665), .C1(new_n501), .C2(new_n502), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n657), .A2(new_n660), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  NOR2_X1   g483(.A1(new_n605), .A2(new_n649), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n642), .A2(new_n503), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  AND2_X1   g486(.A1(new_n503), .A2(new_n438), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n364), .B1(new_n363), .B2(new_n366), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n608), .A2(new_n674), .A3(new_n675), .A4(new_n292), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT104), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G15));
  INV_X1    g494(.A(new_n675), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n291), .A3(new_n367), .A4(new_n607), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n614), .A2(new_n586), .A3(new_n550), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n673), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NOR2_X1   g500(.A1(new_n682), .A2(new_n551), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n641), .A2(new_n586), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n503), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  OAI21_X1  g504(.A(new_n463), .B1(new_n455), .B2(new_n456), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n484), .A2(new_n486), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n488), .B(KEYINPUT105), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n591), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n437), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n674), .A2(new_n675), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n607), .A2(new_n586), .A3(new_n596), .ZN(new_n698));
  INV_X1    g512(.A(new_n550), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n697), .A3(new_n700), .A4(new_n291), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  INV_X1    g516(.A(new_n682), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n641), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT106), .A4(new_n670), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n591), .A2(new_n694), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n670), .A2(new_n631), .A3(new_n634), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n708), .B2(new_n682), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NAND2_X1  g525(.A1(new_n495), .A2(new_n500), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n482), .A2(new_n489), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n438), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n283), .B1(new_n279), .B2(new_n280), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n368), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT42), .A4(new_n670), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n503), .A2(new_n438), .A3(new_n670), .A4(new_n717), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT107), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NAND3_X1  g538(.A1(new_n673), .A2(new_n652), .A3(new_n717), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT108), .B(G134), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G36));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n354), .B2(KEYINPUT45), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n730), .B(new_n344), .C1(new_n349), .C2(new_n353), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT46), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n367), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n360), .B1(new_n351), .B2(new_n352), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n348), .A2(KEYINPUT83), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n337), .A2(new_n343), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n296), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n730), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n354), .A2(KEYINPUT45), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(G469), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT46), .B1(new_n740), .B2(new_n728), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n291), .B(new_n655), .C1(new_n733), .C2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n728), .B1(new_n729), .B2(new_n731), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n367), .A3(new_n732), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT109), .A3(new_n291), .A4(new_n655), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n641), .B2(new_n592), .ZN(new_n752));
  INV_X1    g566(.A(new_n591), .ZN(new_n753));
  INV_X1    g567(.A(new_n498), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n497), .B1(new_n487), .B2(new_n488), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(KEYINPUT110), .A3(new_n631), .A4(new_n634), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n545), .A2(new_n604), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n545), .A2(new_n604), .A3(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n757), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n716), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n716), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n752), .A2(new_n757), .A3(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n750), .A2(new_n765), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  OAI21_X1  g586(.A(new_n291), .B1(new_n733), .B2(new_n741), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n748), .A2(new_n775), .A3(new_n291), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n670), .A2(new_n716), .A3(new_n437), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n503), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  OR3_X1    g594(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT49), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT49), .B1(new_n674), .B2(new_n675), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n758), .A2(new_n292), .A3(new_n283), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n659), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n784), .A2(new_n437), .A3(new_n666), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n697), .A2(new_n291), .A3(new_n716), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n666), .A2(new_n787), .A3(new_n437), .A4(new_n547), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n545), .A2(new_n788), .A3(new_n597), .A4(new_n603), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n762), .A2(new_n646), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n704), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n647), .B1(new_n760), .B2(new_n761), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n659), .A2(new_n793), .A3(new_n283), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n696), .A2(new_n291), .A3(new_n697), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n793), .A2(new_n696), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n716), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n774), .A2(new_n776), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n674), .A2(new_n675), .A3(new_n291), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT113), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n786), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n789), .A2(new_n799), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n804), .B1(new_n774), .B2(new_n776), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n808), .B(KEYINPUT51), .C1(new_n802), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n791), .A2(new_n715), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT114), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n791), .A2(new_n813), .A3(new_n715), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n801), .A2(new_n703), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(G952), .A3(new_n187), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n788), .B2(new_n606), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(KEYINPUT48), .A3(new_n814), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n807), .B(new_n810), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n701), .B1(new_n369), .B2(new_n635), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n605), .B1(new_n585), .B2(new_n596), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n438), .A3(new_n592), .A4(new_n550), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n369), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n438), .B(new_n503), .C1(new_n676), .C2(new_n684), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n689), .A4(new_n588), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n503), .A2(new_n688), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n708), .B1(new_n836), .B2(new_n651), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n717), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n710), .A2(new_n653), .A3(new_n671), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n434), .A2(new_n633), .A3(new_n650), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n698), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n666), .A2(new_n368), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n723), .A2(new_n725), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n844), .B(KEYINPUT112), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n851), .B2(new_n839), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n838), .A2(new_n852), .A3(new_n847), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(new_n849), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n853), .B2(new_n857), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n827), .A2(new_n828), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n785), .B1(new_n860), .B2(new_n861), .ZN(G75));
  AOI21_X1  g676(.A(new_n366), .B1(new_n853), .B2(new_n857), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n276), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n268), .A2(new_n272), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n270), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n187), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G51));
  XOR2_X1   g686(.A(new_n728), .B(KEYINPUT57), .Z(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n858), .B2(new_n859), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n363), .ZN(new_n875));
  INV_X1    g689(.A(new_n863), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(new_n740), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n871), .B1(new_n875), .B2(new_n877), .ZN(G54));
  AND2_X1   g692(.A1(new_n532), .A2(new_n540), .ZN(new_n879));
  NAND2_X1  g693(.A1(KEYINPUT58), .A2(G475), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n863), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n863), .B2(new_n881), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n871), .ZN(G60));
  NAND2_X1  g698(.A1(G478), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n858), .B2(new_n859), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n600), .A2(new_n602), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n871), .ZN(new_n890));
  INV_X1    g704(.A(new_n888), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n886), .C1(new_n858), .C2(new_n859), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(G63));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT60), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n853), .B2(new_n857), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n628), .B(KEYINPUT117), .Z(new_n897));
  AOI21_X1  g711(.A(new_n871), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT118), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  OAI221_X1 g713(.A(new_n898), .B1(new_n430), .B2(new_n896), .C1(new_n899), .C2(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n897), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n901), .B(new_n890), .C1(new_n430), .C2(new_n896), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT61), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(G66));
  AOI21_X1  g720(.A(new_n187), .B1(new_n549), .B2(G224), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n835), .B(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n910), .B2(new_n187), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n866), .B1(G898), .B2(new_n187), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n911), .B(new_n912), .Z(G69));
  NAND2_X1  g727(.A1(new_n471), .A2(new_n472), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(new_n536), .Z(new_n915));
  INV_X1    g729(.A(G900), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n187), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n771), .A2(new_n918), .A3(new_n840), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n771), .B2(new_n840), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n774), .A2(new_n778), .A3(new_n776), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n714), .A2(new_n698), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n744), .B2(new_n749), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n925), .A2(new_n723), .A3(new_n725), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n927), .B2(new_n187), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n668), .A2(new_n710), .A3(new_n653), .A4(new_n671), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  INV_X1    g744(.A(new_n656), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n673), .A2(new_n931), .A3(new_n716), .A4(new_n830), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n932), .A2(new_n779), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n771), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT120), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n929), .B(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n771), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n915), .B1(new_n940), .B2(new_n187), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n928), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n294), .B2(new_n916), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n915), .B2(KEYINPUT122), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n942), .B(new_n945), .ZN(G72));
  NAND2_X1  g760(.A1(G472), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  XOR2_X1   g762(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n940), .B2(new_n910), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n853), .A2(new_n857), .ZN(new_n952));
  INV_X1    g766(.A(new_n661), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n474), .A2(new_n463), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n950), .ZN(new_n955));
  AOI22_X1  g769(.A1(new_n951), .A2(new_n661), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(KEYINPUT126), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n926), .B(new_n909), .C1(new_n920), .C2(new_n919), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n950), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n961), .A3(new_n950), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n871), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g779(.A(KEYINPUT127), .B(new_n871), .C1(new_n960), .C2(new_n962), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G57));
endmodule


