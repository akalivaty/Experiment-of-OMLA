//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G952), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  INV_X1    g005(.A(G234), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT21), .B(G898), .Z(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(KEYINPUT96), .ZN(new_n197));
  INV_X1    g011(.A(G902), .ZN(new_n198));
  INV_X1    g012(.A(G953), .ZN(new_n199));
  AOI211_X1 g013(.A(new_n198), .B(new_n199), .C1(G234), .C2(G237), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n195), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G214), .B1(G237), .B2(G902), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(G116), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT2), .A2(G113), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT2), .A2(G113), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n218), .B(new_n219), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(G116), .A2(G119), .ZN(new_n227));
  NOR2_X1   g041(.A1(G116), .A2(G119), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n226), .B(new_n220), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n211), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n216), .A2(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G113), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n227), .A2(new_n228), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n234), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT87), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n225), .B1(new_n234), .B2(new_n235), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n241), .B(new_n242), .C1(new_n238), .C2(new_n234), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n229), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n208), .A2(G104), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n205), .A2(G107), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n214), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT81), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n214), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n233), .B1(new_n244), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G122), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n233), .C1(new_n244), .C2(new_n252), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(KEYINPUT6), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT0), .B(G128), .Z(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n264), .B(G125), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n261), .B(G146), .C1(new_n268), .C2(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n259), .A3(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n268), .A2(KEYINPUT1), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n260), .A3(new_n262), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n267), .B1(new_n275), .B2(G125), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n199), .A2(G224), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n253), .A2(new_n279), .A3(new_n255), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n258), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n267), .B2(KEYINPUT88), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  OAI221_X1 g098(.A(new_n267), .B1(KEYINPUT88), .B2(new_n282), .C1(new_n275), .C2(G125), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n214), .A2(new_n247), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n244), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n254), .B(KEYINPUT8), .Z(new_n289));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n238), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n229), .B1(new_n237), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n286), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n294), .B2(new_n257), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n281), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n296), .B(KEYINPUT89), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n281), .B2(new_n295), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n204), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n198), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n273), .A2(new_n260), .A3(new_n262), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT66), .B1(new_n305), .B2(new_n271), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n274), .A2(new_n307), .A3(new_n269), .A4(new_n270), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n306), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n214), .A2(new_n247), .A3(new_n250), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n250), .B1(new_n214), .B2(new_n247), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n211), .A2(G101), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n314), .B(new_n232), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT11), .B1(new_n318), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G134), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT64), .B1(new_n321), .B2(G134), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT64), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n318), .A3(G137), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n323), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT82), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n266), .A2(new_n339), .A3(new_n273), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n272), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n287), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n313), .A2(new_n317), .A3(new_n337), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT83), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n232), .A2(new_n314), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n343), .A2(new_n342), .B1(new_n347), .B2(new_n215), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n313), .A4(new_n337), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n199), .A2(G227), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(G140), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT79), .B(G110), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n348), .A2(new_n313), .B1(new_n335), .B2(new_n333), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n333), .A2(new_n335), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n271), .B1(KEYINPUT80), .B2(new_n274), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n248), .B1(new_n361), .B2(new_n340), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n287), .A2(new_n275), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT12), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n317), .B1(new_n362), .B2(KEYINPUT10), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n306), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n252), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n349), .B1(new_n370), .B2(new_n337), .ZN(new_n371));
  INV_X1    g185(.A(new_n350), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n355), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n364), .B(KEYINPUT12), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n350), .B2(new_n346), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT84), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n359), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n304), .B1(new_n379), .B2(G469), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n351), .A2(new_n357), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n382));
  INV_X1    g196(.A(new_n355), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n351), .A2(new_n355), .A3(new_n366), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n356), .B1(new_n346), .B2(new_n350), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT85), .B1(new_n386), .B2(new_n355), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n303), .A3(new_n198), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n189), .B(new_n302), .C1(new_n380), .C2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G472), .A2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n318), .A2(G137), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n321), .A2(G134), .ZN(new_n394));
  OAI21_X1  g208(.A(G131), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n306), .A2(new_n335), .A3(new_n395), .A4(new_n308), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n314), .B1(new_n329), .B2(new_n330), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n223), .A2(new_n229), .A3(KEYINPUT67), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT67), .B1(new_n223), .B2(new_n229), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(G237), .A2(G953), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT27), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G210), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n402), .B2(G210), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT26), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT26), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n407), .A2(new_n410), .A3(G101), .ZN(new_n411));
  AOI21_X1  g225(.A(G101), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n335), .A2(new_n395), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT65), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n335), .A2(KEYINPUT65), .A3(new_n395), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n275), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT30), .B1(new_n420), .B2(new_n397), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n230), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n414), .B(new_n415), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(KEYINPUT0), .A2(G128), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n260), .A2(new_n262), .B1(new_n426), .B2(new_n263), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n333), .B2(new_n335), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n305), .A2(new_n271), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n416), .B2(new_n417), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n432), .B2(new_n419), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n230), .B(new_n422), .C1(new_n433), .C2(KEYINPUT30), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n415), .B1(new_n434), .B2(new_n414), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT31), .B1(new_n425), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n414), .B1(new_n421), .B2(new_n423), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT31), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n441));
  AOI22_X1  g255(.A1(new_n420), .A2(new_n397), .B1(new_n223), .B2(new_n229), .ZN(new_n442));
  INV_X1    g256(.A(new_n401), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(KEYINPUT28), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n413), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n392), .B1(new_n440), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n446), .A3(new_n413), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT71), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n444), .A2(new_n446), .A3(new_n453), .A4(new_n413), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n434), .A2(new_n401), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT72), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n401), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n397), .A2(new_n396), .A3(new_n400), .A4(KEYINPUT72), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n396), .A2(new_n397), .ZN(new_n462));
  INV_X1    g276(.A(new_n400), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT73), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT73), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n445), .B1(new_n468), .B2(KEYINPUT28), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n413), .A2(KEYINPUT29), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n450), .A2(KEYINPUT32), .B1(new_n472), .B2(G472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT70), .B1(new_n450), .B2(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n437), .A2(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n438), .B1(new_n475), .B2(new_n424), .ZN(new_n476));
  INV_X1    g290(.A(new_n439), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n449), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n391), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT23), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n217), .B2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n217), .A2(G128), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n268), .A2(KEYINPUT23), .A3(G119), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G110), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT75), .B1(new_n217), .B2(G128), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT75), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n268), .A3(G119), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n494), .A3(new_n487), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT24), .B(G110), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n490), .A2(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT77), .A2(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G140), .ZN(new_n499));
  INV_X1    g313(.A(G140), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT77), .A3(G125), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT16), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT16), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n500), .A3(G125), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(G146), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G125), .B(G140), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n259), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n484), .B1(new_n497), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n495), .A2(new_n496), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(G110), .B2(new_n489), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n511), .A2(KEYINPUT78), .A3(new_n505), .A4(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n502), .A2(new_n504), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n259), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n505), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n491), .B1(new_n489), .B2(KEYINPUT76), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(KEYINPUT76), .B2(new_n489), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n518), .C1(new_n496), .C2(new_n495), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT22), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(G137), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n519), .A3(new_n523), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n198), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT25), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n529), .A3(new_n198), .A4(new_n526), .ZN(new_n530));
  OAI21_X1  g344(.A(G217), .B1(new_n192), .B2(G902), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n525), .A2(new_n526), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n532), .A2(G902), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n205), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n499), .A2(new_n501), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n507), .B1(new_n542), .B2(new_n259), .ZN(new_n543));
  AND4_X1   g357(.A1(G143), .A2(new_n193), .A3(new_n199), .A4(G214), .ZN(new_n544));
  AOI21_X1  g358(.A(G143), .B1(new_n402), .B2(G214), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT18), .B(G131), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n193), .A2(new_n199), .A3(G214), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n261), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n402), .A2(G143), .A3(G214), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT18), .A2(G131), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT17), .B(G131), .C1(new_n544), .C2(new_n545), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n515), .A2(new_n505), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G131), .B1(new_n544), .B2(new_n545), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n328), .A3(new_n549), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n541), .B(new_n552), .C1(new_n554), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(new_n505), .A3(new_n515), .A4(new_n553), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT90), .A3(new_n541), .A4(new_n552), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n555), .A2(new_n557), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n506), .A2(KEYINPUT19), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(KEYINPUT19), .B2(new_n542), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n505), .B(new_n566), .C1(new_n568), .C2(G146), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n552), .ZN(new_n570));
  INV_X1    g384(.A(new_n541), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n574));
  NOR2_X1   g388(.A1(G475), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n575), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT20), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n541), .B1(new_n563), .B2(new_n552), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n561), .B2(new_n564), .ZN(new_n583));
  OAI21_X1  g397(.A(G475), .B1(new_n583), .B2(G902), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n187), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(G217), .A3(new_n199), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n216), .B2(G122), .ZN(new_n589));
  INV_X1    g403(.A(G122), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT92), .A3(G116), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n216), .A2(G122), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n592), .A2(new_n208), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n208), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g410(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n597), .A2(G128), .A3(new_n261), .A4(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n600));
  NAND2_X1  g414(.A1(new_n268), .A2(G143), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n261), .A2(G128), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n599), .B(G134), .C1(new_n600), .C2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n318), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(G134), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n605), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n592), .A2(new_n208), .A3(new_n593), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT14), .B1(new_n590), .B2(G116), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT14), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n216), .A3(G122), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n592), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT94), .A3(G107), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT94), .B1(new_n616), .B2(G107), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n607), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n589), .A2(new_n591), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n613), .A2(new_n615), .ZN(new_n624));
  OAI21_X1  g438(.A(G107), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n611), .B1(new_n627), .B2(new_n617), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n596), .A2(new_n606), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT95), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n587), .B1(new_n622), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n587), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n621), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n198), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT15), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n585), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n390), .A2(new_n483), .A3(new_n539), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  NAND2_X1  g455(.A1(new_n281), .A2(new_n295), .ZN(new_n642));
  INV_X1    g456(.A(new_n296), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n203), .B1(new_n644), .B2(new_n297), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n636), .A2(G902), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n631), .A2(new_n634), .A3(KEYINPUT33), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n632), .B1(new_n633), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(KEYINPUT97), .B(new_n587), .C1(new_n628), .C2(new_n629), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n647), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n635), .A2(new_n636), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n585), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n646), .A2(new_n657), .A3(new_n201), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n189), .B1(new_n380), .B2(new_n389), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n478), .B2(new_n198), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n661), .A2(new_n450), .A3(new_n538), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n578), .A2(new_n584), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n574), .A2(new_n577), .ZN(new_n668));
  INV_X1    g482(.A(new_n575), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n580), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n638), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n666), .B1(new_n671), .B2(new_n201), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n670), .A2(new_n578), .A3(new_n584), .ZN(new_n673));
  INV_X1    g487(.A(new_n201), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(KEYINPUT98), .A3(new_n638), .A4(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n672), .A2(new_n675), .A3(new_n645), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n659), .A3(new_n662), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n524), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n520), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n536), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n533), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n533), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n661), .A3(new_n450), .ZN(new_n688));
  INV_X1    g502(.A(new_n204), .ZN(new_n689));
  INV_X1    g503(.A(new_n301), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(new_n297), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n659), .A3(new_n639), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AOI21_X1  g508(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n695));
  AOI211_X1 g509(.A(KEYINPUT70), .B(KEYINPUT32), .C1(new_n478), .C2(new_n391), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n687), .B1(new_n697), .B2(new_n473), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n195), .B1(new_n200), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n671), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n659), .A2(new_n645), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(new_n700), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n659), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n468), .A2(new_n448), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n475), .A3(new_n424), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n660), .B1(new_n709), .B2(new_n198), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n450), .B2(KEYINPUT32), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n697), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n585), .A2(new_n638), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n690), .A2(new_n297), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n533), .A3(new_n202), .A4(new_n682), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n707), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  INV_X1    g534(.A(new_n700), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n585), .A2(new_n656), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n585), .A2(new_n656), .A3(KEYINPUT100), .A4(new_n721), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n698), .A2(new_n702), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  AOI21_X1  g542(.A(new_n538), .B1(new_n697), .B2(new_n473), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n388), .A2(new_n198), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT101), .A3(new_n389), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n733), .A3(G469), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n189), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n729), .A2(new_n658), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n736), .B(new_n738), .ZN(G15));
  NAND3_X1  g553(.A1(new_n729), .A2(new_n676), .A3(new_n735), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n645), .ZN(new_n742));
  INV_X1    g556(.A(new_n687), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n483), .A2(new_n639), .A3(new_n674), .A4(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND2_X1  g560(.A1(new_n732), .A2(new_n734), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n475), .A2(new_n424), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n477), .B1(new_n748), .B2(KEYINPUT31), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n469), .A2(new_n413), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n391), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(G902), .B1(new_n440), .B2(new_n449), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n539), .B(new_n751), .C1(new_n752), .C2(new_n660), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n645), .A2(new_n638), .A3(new_n585), .A4(new_n674), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n747), .A2(new_n755), .A3(new_n188), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  INV_X1    g571(.A(new_n661), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n683), .A3(new_n751), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n724), .A2(new_n725), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n735), .A3(new_n645), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NAND4_X1  g577(.A1(new_n690), .A2(new_n188), .A3(new_n297), .A4(new_n202), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n538), .B(new_n764), .C1(new_n380), .C2(new_n389), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n726), .A3(new_n483), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT103), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n479), .A2(new_n771), .A3(new_n481), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT104), .B1(new_n450), .B2(KEYINPUT32), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n473), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n539), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n380), .A2(new_n389), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n777), .A2(new_n768), .A3(new_n764), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n726), .ZN(new_n779));
  OAI22_X1  g593(.A1(new_n769), .A2(new_n770), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  AND2_X1   g595(.A1(new_n765), .A2(new_n483), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n701), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  OAI21_X1  g598(.A(new_n383), .B1(new_n377), .B2(KEYINPUT84), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n373), .A2(new_n374), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n358), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n379), .A2(KEYINPUT45), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(G469), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n303), .B2(new_n198), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n389), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n188), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n656), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n585), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(KEYINPUT105), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n758), .A2(new_n479), .B1(new_n533), .B2(new_n682), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT44), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n690), .A2(new_n297), .A3(new_n202), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT106), .Z(new_n811));
  NAND4_X1  g625(.A1(new_n798), .A2(new_n809), .A3(new_n705), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  XNOR2_X1  g627(.A(new_n797), .B(KEYINPUT47), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n483), .A2(new_n539), .A3(new_n810), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n726), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n810), .A2(new_n638), .A3(new_n700), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n698), .A2(new_n659), .A3(new_n673), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n777), .A2(new_n764), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n761), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n783), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n780), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n657), .B(KEYINPUT107), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n390), .A2(new_n662), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n640), .A2(new_n756), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n667), .A2(new_n638), .A3(new_n581), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n302), .ZN(new_n832));
  INV_X1    g646(.A(new_n585), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n691), .A2(KEYINPUT108), .A3(new_n833), .A4(new_n638), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n659), .A2(new_n832), .A3(new_n662), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n829), .B1(new_n692), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n729), .B(new_n735), .C1(new_n676), .C2(new_n658), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n692), .A2(new_n835), .A3(new_n829), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n745), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n819), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n783), .A2(new_n821), .A3(new_n823), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n766), .A2(new_n768), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT103), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n779), .A2(new_n775), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n692), .A2(new_n835), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT109), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n639), .A2(new_n776), .A3(new_n188), .A4(new_n691), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n729), .A2(new_n851), .B1(new_n735), .B2(new_n755), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n852), .A3(new_n839), .A4(new_n827), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n838), .B1(new_n742), .B2(new_n744), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n855), .A3(KEYINPUT110), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n857), .B2(KEYINPUT111), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n841), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n698), .B(new_n702), .C1(new_n701), .C2(new_n726), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n646), .A2(new_n714), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n683), .A2(new_n700), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n659), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n865), .B2(new_n712), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n762), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n861), .A2(new_n866), .A3(KEYINPUT112), .A4(new_n762), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n712), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n861), .A2(new_n762), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(KEYINPUT114), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n858), .A2(new_n860), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n862), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n867), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n841), .A2(new_n856), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT53), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n825), .A2(new_n840), .A3(new_n887), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n871), .A2(KEYINPUT114), .A3(new_n875), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT114), .B1(new_n871), .B2(new_n875), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n735), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n810), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n194), .B1(new_n803), .B2(new_n805), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n775), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT48), .ZN(new_n900));
  INV_X1    g714(.A(new_n753), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n712), .A2(new_n538), .A3(new_n194), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  OAI221_X1 g718(.A(new_n191), .B1(new_n742), .B2(new_n902), .C1(new_n904), .C2(new_n657), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n898), .A2(new_n759), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n896), .A2(new_n903), .A3(new_n833), .A4(new_n799), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n895), .A2(new_n202), .A3(new_n716), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(KEYINPUT50), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n909), .A2(new_n902), .A3(new_n912), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n907), .B(new_n908), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n897), .A2(new_n901), .A3(new_n811), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n747), .A2(new_n189), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n814), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n906), .B1(new_n920), .B2(KEYINPUT51), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n907), .A2(new_n908), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(KEYINPUT51), .C1(new_n915), .C2(new_n914), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n814), .A2(new_n918), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n924), .B2(KEYINPUT116), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n886), .A2(new_n894), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT117), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n886), .A2(new_n928), .A3(new_n931), .A4(new_n894), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n190), .A2(new_n199), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT49), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n747), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n732), .A2(KEYINPUT49), .A3(new_n734), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n539), .A2(new_n188), .A3(new_n202), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n716), .A2(new_n801), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n713), .A2(new_n936), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(new_n940), .ZN(G75));
  NOR2_X1   g755(.A1(new_n199), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n888), .A2(new_n892), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(G902), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n300), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n258), .A2(new_n280), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(new_n278), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT56), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(G210), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n945), .A2(KEYINPUT118), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT118), .B1(new_n945), .B2(new_n952), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n956), .B2(new_n949), .ZN(G51));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n880), .A2(new_n889), .B1(new_n884), .B2(new_n887), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n959), .A2(new_n198), .A3(new_n791), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n304), .B(KEYINPUT57), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n888), .A2(new_n892), .A3(new_n893), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n893), .B1(new_n888), .B2(new_n892), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n964), .B2(new_n388), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n958), .B1(new_n965), .B2(new_n942), .ZN(new_n966));
  INV_X1    g780(.A(new_n388), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n894), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n961), .ZN(new_n970));
  OAI211_X1 g784(.A(KEYINPUT119), .B(new_n943), .C1(new_n970), .C2(new_n960), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n966), .A2(new_n971), .ZN(G54));
  NAND2_X1  g786(.A1(KEYINPUT58), .A2(G475), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT120), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n944), .A2(G902), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n943), .B1(new_n975), .B2(new_n668), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n668), .B2(new_n975), .ZN(G60));
  OR2_X1    g791(.A1(new_n648), .A2(new_n653), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n886), .A2(new_n894), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT59), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n969), .A2(new_n978), .A3(new_n981), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n942), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n888), .B2(new_n892), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT121), .B1(new_n987), .B2(new_n681), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(KEYINPUT61), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n942), .B1(new_n987), .B2(new_n681), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT122), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n534), .B1(new_n959), .B2(new_n986), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n986), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n944), .A2(new_n681), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n943), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n987), .A2(new_n535), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT122), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1001), .A2(new_n989), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n996), .A2(new_n1003), .ZN(G66));
  NOR2_X1   g818(.A1(new_n855), .A2(G953), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  INV_X1    g820(.A(G224), .ZN(new_n1007));
  OAI21_X1  g821(.A(G953), .B1(new_n197), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n947), .B1(G898), .B2(new_n199), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  INV_X1    g825(.A(new_n719), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n861), .A2(new_n762), .ZN(new_n1013));
  OR3_X1    g827(.A1(new_n1012), .A2(KEYINPUT62), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT62), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  INV_X1    g829(.A(new_n831), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n782), .B(new_n705), .C1(new_n1016), .C2(new_n826), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n812), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n817), .A2(new_n1014), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n199), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n422), .B1(new_n433), .B2(KEYINPUT30), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT124), .Z(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT125), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(new_n568), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(G900), .B2(G953), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n812), .A2(new_n783), .ZN(new_n1027));
  INV_X1    g841(.A(new_n775), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n705), .A2(new_n798), .A3(new_n863), .A4(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1029), .A2(new_n1013), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n817), .A2(new_n780), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1026), .B1(new_n1031), .B2(G953), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n199), .B1(G227), .B2(G900), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1034), .B1(new_n1032), .B2(KEYINPUT126), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1033), .B(new_n1035), .Z(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n1031), .B2(new_n840), .ZN(new_n1039));
  INV_X1    g853(.A(new_n455), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1039), .A2(new_n448), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1038), .B1(new_n1019), .B2(new_n840), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1042), .A2(new_n413), .A3(new_n455), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1041), .A2(new_n1043), .A3(new_n943), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n881), .A2(new_n885), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1038), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1040), .A2(new_n413), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  OR2_X1    g862(.A1(new_n1048), .A2(KEYINPUT127), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n748), .B1(new_n1048), .B2(KEYINPUT127), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1044), .B1(new_n1045), .B2(new_n1051), .ZN(G57));
endmodule


