

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n358, n359, n360, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n485, n486, n487,
         n488, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769;

  AND2_X1 U373 ( .A1(n352), .A2(n351), .ZN(n610) );
  INV_X1 U374 ( .A(n608), .ZN(n351) );
  INV_X1 U375 ( .A(n597), .ZN(n353) );
  INV_X1 U376 ( .A(KEYINPUT34), .ZN(n354) );
  XNOR2_X1 U377 ( .A(n410), .B(n463), .ZN(n648) );
  XNOR2_X1 U378 ( .A(n504), .B(n506), .ZN(n392) );
  XNOR2_X1 U379 ( .A(n569), .B(KEYINPUT75), .ZN(n369) );
  NAND2_X2 U380 ( .A1(n380), .A2(n595), .ZN(n598) );
  XNOR2_X1 U381 ( .A(n598), .B(n353), .ZN(n352) );
  AND2_X2 U382 ( .A1(n404), .A2(n412), .ZN(n411) );
  XNOR2_X2 U383 ( .A(n596), .B(KEYINPUT73), .ZN(n597) );
  NOR2_X2 U384 ( .A1(n702), .A2(n701), .ZN(n572) );
  XNOR2_X1 U385 ( .A(n625), .B(KEYINPUT76), .ZN(n440) );
  NOR2_X2 U386 ( .A1(n377), .A2(n402), .ZN(n599) );
  AND2_X2 U387 ( .A1(n748), .A2(n628), .ZN(n629) );
  NOR2_X2 U388 ( .A1(n600), .A2(n611), .ZN(n601) );
  XNOR2_X1 U389 ( .A(n355), .B(n354), .ZN(n433) );
  NAND2_X1 U390 ( .A1(n373), .A2(n380), .ZN(n355) );
  XNOR2_X2 U391 ( .A(n356), .B(KEYINPUT65), .ZN(n647) );
  NAND2_X2 U392 ( .A1(n446), .A2(n447), .ZN(n356) );
  XNOR2_X2 U393 ( .A(n557), .B(n556), .ZN(n574) );
  XNOR2_X1 U394 ( .A(n358), .B(n485), .ZN(n416) );
  XNOR2_X1 U395 ( .A(n483), .B(n521), .ZN(n358) );
  XNOR2_X2 U396 ( .A(n359), .B(n375), .ZN(n581) );
  NAND2_X1 U397 ( .A1(n396), .A2(n427), .ZN(n359) );
  XNOR2_X2 U398 ( .A(n360), .B(n488), .ZN(n709) );
  NAND2_X2 U399 ( .A1(n415), .A2(n496), .ZN(n360) );
  XNOR2_X2 U400 ( .A(KEYINPUT24), .B(G137), .ZN(n480) );
  XNOR2_X2 U401 ( .A(n436), .B(n435), .ZN(n643) );
  NOR2_X2 U402 ( .A1(n578), .A2(n378), .ZN(n549) );
  XNOR2_X2 U403 ( .A(n543), .B(n544), .ZN(n611) );
  INV_X1 U404 ( .A(n647), .ZN(n667) );
  XOR2_X1 U405 ( .A(KEYINPUT97), .B(KEYINPUT94), .Z(n515) );
  INV_X2 U406 ( .A(G953), .ZN(n758) );
  BUF_X1 U407 ( .A(G122), .Z(n528) );
  NOR2_X2 U408 ( .A1(n566), .A2(n565), .ZN(n370) );
  OR2_X2 U409 ( .A1(n648), .A2(G902), .ZN(n464) );
  AND2_X2 U410 ( .A1(n538), .A2(n558), .ZN(n688) );
  NOR2_X2 U411 ( .A1(G902), .A2(n633), .ZN(n525) );
  INV_X4 U412 ( .A(G143), .ZN(n454) );
  XNOR2_X1 U413 ( .A(n437), .B(KEYINPUT42), .ZN(n769) );
  XNOR2_X1 U414 ( .A(G119), .B(KEYINPUT23), .ZN(n477) );
  INV_X1 U415 ( .A(KEYINPUT76), .ZN(n363) );
  AND2_X1 U416 ( .A1(n629), .A2(n631), .ZN(n448) );
  XNOR2_X1 U417 ( .A(n366), .B(KEYINPUT46), .ZN(n365) );
  NOR2_X2 U418 ( .A1(n643), .A2(n769), .ZN(n366) );
  NOR2_X1 U419 ( .A1(n473), .A2(n428), .ZN(n385) );
  BUF_X1 U420 ( .A(n615), .Z(n402) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X1 U422 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n501) );
  XNOR2_X1 U423 ( .A(G110), .B(G128), .ZN(n478) );
  INV_X2 U424 ( .A(KEYINPUT67), .ZN(n407) );
  XNOR2_X1 U425 ( .A(n627), .B(n363), .ZN(n364) );
  XNOR2_X2 U426 ( .A(n586), .B(KEYINPUT81), .ZN(n627) );
  NAND2_X1 U427 ( .A1(n364), .A2(n448), .ZN(n447) );
  NAND2_X1 U428 ( .A1(n364), .A2(n629), .ZN(n735) );
  NAND2_X2 U429 ( .A1(n367), .A2(n365), .ZN(n371) );
  XNOR2_X2 U430 ( .A(n368), .B(KEYINPUT69), .ZN(n367) );
  NAND2_X1 U431 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X2 U432 ( .A(n371), .B(n398), .ZN(n394) );
  INV_X1 U433 ( .A(n380), .ZN(n376) );
  XNOR2_X2 U434 ( .A(n592), .B(n372), .ZN(n380) );
  INV_X1 U435 ( .A(KEYINPUT0), .ZN(n372) );
  INV_X1 U436 ( .A(n697), .ZN(n373) );
  AND2_X1 U437 ( .A1(n767), .A2(n444), .ZN(n443) );
  INV_X1 U438 ( .A(KEYINPUT48), .ZN(n398) );
  XNOR2_X1 U439 ( .A(KEYINPUT15), .B(G902), .ZN(n630) );
  XNOR2_X1 U440 ( .A(n504), .B(G137), .ZN(n434) );
  XNOR2_X1 U441 ( .A(n474), .B(KEYINPUT8), .ZN(n526) );
  NOR2_X1 U442 ( .A1(n417), .A2(G953), .ZN(n474) );
  INV_X1 U443 ( .A(G234), .ZN(n417) );
  XNOR2_X1 U444 ( .A(n430), .B(G107), .ZN(n529) );
  INV_X1 U445 ( .A(G116), .ZN(n430) );
  INV_X1 U446 ( .A(KEYINPUT2), .ZN(n439) );
  INV_X1 U447 ( .A(n416), .ZN(n415) );
  INV_X1 U448 ( .A(KEYINPUT93), .ZN(n458) );
  XOR2_X1 U449 ( .A(KEYINPUT5), .B(G131), .Z(n457) );
  XNOR2_X1 U450 ( .A(G113), .B(G116), .ZN(n456) );
  XOR2_X1 U451 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n527) );
  INV_X1 U452 ( .A(KEYINPUT100), .ZN(n423) );
  NAND2_X1 U453 ( .A1(n526), .A2(G217), .ZN(n424) );
  XNOR2_X1 U454 ( .A(n453), .B(n518), .ZN(n519) );
  XNOR2_X1 U455 ( .A(n572), .B(n571), .ZN(n730) );
  XNOR2_X1 U456 ( .A(n465), .B(KEYINPUT30), .ZN(n473) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X1 U458 ( .A(n432), .B(n431), .ZN(n444) );
  INV_X1 U459 ( .A(KEYINPUT35), .ZN(n431) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n466) );
  OR2_X1 U461 ( .A1(G237), .A2(G902), .ZN(n507) );
  INV_X1 U462 ( .A(KEYINPUT44), .ZN(n441) );
  AND2_X1 U463 ( .A1(n626), .A2(KEYINPUT2), .ZN(n449) );
  XOR2_X1 U464 ( .A(n515), .B(n514), .Z(n453) );
  XNOR2_X1 U465 ( .A(KEYINPUT98), .B(KEYINPUT11), .ZN(n514) );
  XNOR2_X1 U466 ( .A(G143), .B(G104), .ZN(n516) );
  XOR2_X1 U467 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n517) );
  XOR2_X1 U468 ( .A(G131), .B(G140), .Z(n522) );
  XNOR2_X1 U469 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n758), .A2(G224), .ZN(n405) );
  AND2_X1 U471 ( .A1(n414), .A2(n699), .ZN(n396) );
  XNOR2_X1 U472 ( .A(n573), .B(n550), .ZN(n615) );
  INV_X1 U473 ( .A(KEYINPUT1), .ZN(n550) );
  INV_X1 U474 ( .A(KEYINPUT22), .ZN(n596) );
  INV_X1 U475 ( .A(n585), .ZN(n397) );
  BUF_X1 U476 ( .A(n697), .Z(n731) );
  XNOR2_X1 U477 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n475) );
  XNOR2_X1 U478 ( .A(n424), .B(n422), .ZN(n534) );
  XNOR2_X1 U479 ( .A(n527), .B(n423), .ZN(n422) );
  AND2_X1 U480 ( .A1(n419), .A2(n418), .ZN(n696) );
  XNOR2_X1 U481 ( .A(n420), .B(KEYINPUT43), .ZN(n419) );
  NOR2_X1 U482 ( .A1(n730), .A2(n575), .ZN(n437) );
  INV_X1 U483 ( .A(KEYINPUT40), .ZN(n435) );
  XNOR2_X1 U484 ( .A(n384), .B(KEYINPUT105), .ZN(n383) );
  NAND2_X1 U485 ( .A1(n385), .A2(n414), .ZN(n384) );
  INV_X1 U486 ( .A(n574), .ZN(n413) );
  INV_X1 U487 ( .A(KEYINPUT60), .ZN(n450) );
  INV_X1 U488 ( .A(n444), .ZN(n765) );
  AND2_X1 U489 ( .A1(n620), .A2(n709), .ZN(n374) );
  INV_X1 U490 ( .A(G902), .ZN(n496) );
  XNOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n375) );
  NOR2_X1 U492 ( .A1(n473), .A2(n472), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n598), .B(n597), .ZN(n377) );
  BUF_X1 U494 ( .A(n554), .Z(n378) );
  BUF_X1 U495 ( .A(n748), .Z(n379) );
  INV_X1 U496 ( .A(n376), .ZN(n618) );
  INV_X1 U497 ( .A(n547), .ZN(n580) );
  XNOR2_X1 U498 ( .A(n580), .B(KEYINPUT38), .ZN(n576) );
  NAND2_X1 U499 ( .A1(n580), .A2(n539), .ZN(n428) );
  XNOR2_X1 U500 ( .A(n741), .B(n386), .ZN(n381) );
  XNOR2_X1 U501 ( .A(n741), .B(n386), .ZN(n656) );
  XNOR2_X2 U502 ( .A(n382), .B(G134), .ZN(n530) );
  XNOR2_X1 U503 ( .A(n390), .B(n382), .ZN(n389) );
  XNOR2_X2 U504 ( .A(n454), .B(G128), .ZN(n382) );
  NAND2_X1 U505 ( .A1(n383), .A2(n603), .ZN(n646) );
  XNOR2_X2 U506 ( .A(n387), .B(n389), .ZN(n386) );
  XNOR2_X2 U507 ( .A(n392), .B(n391), .ZN(n387) );
  XNOR2_X2 U508 ( .A(n388), .B(n503), .ZN(n741) );
  XNOR2_X2 U509 ( .A(n393), .B(n529), .ZN(n388) );
  XNOR2_X1 U510 ( .A(n406), .B(KEYINPUT18), .ZN(n390) );
  XNOR2_X2 U511 ( .A(n505), .B(n405), .ZN(n391) );
  XNOR2_X2 U512 ( .A(n500), .B(n501), .ZN(n393) );
  AND2_X1 U513 ( .A1(n394), .A2(n397), .ZN(n628) );
  NAND2_X1 U514 ( .A1(n394), .A2(n438), .ZN(n586) );
  NAND2_X1 U515 ( .A1(n581), .A2(n688), .ZN(n436) );
  XNOR2_X1 U516 ( .A(n610), .B(n609), .ZN(n767) );
  INV_X2 U517 ( .A(KEYINPUT3), .ZN(n429) );
  XNOR2_X1 U518 ( .A(n442), .B(n441), .ZN(n400) );
  XNOR2_X2 U519 ( .A(n399), .B(KEYINPUT77), .ZN(n639) );
  NAND2_X1 U520 ( .A1(n411), .A2(n413), .ZN(n399) );
  NAND2_X1 U521 ( .A1(n400), .A2(n624), .ZN(n409) );
  XNOR2_X1 U522 ( .A(n401), .B(n753), .ZN(n633) );
  XNOR2_X1 U523 ( .A(n519), .B(n520), .ZN(n401) );
  NAND2_X1 U524 ( .A1(n694), .A2(n552), .ZN(n566) );
  NAND2_X1 U525 ( .A1(n551), .A2(n607), .ZN(n694) );
  XNOR2_X2 U526 ( .A(n525), .B(n524), .ZN(n538) );
  NAND2_X1 U527 ( .A1(n443), .A2(n645), .ZN(n442) );
  INV_X2 U528 ( .A(KEYINPUT4), .ZN(n408) );
  NOR2_X1 U529 ( .A1(n711), .A2(n573), .ZN(n403) );
  NAND2_X1 U530 ( .A1(n404), .A2(n591), .ZN(n592) );
  XNOR2_X1 U531 ( .A(n554), .B(n553), .ZN(n404) );
  XNOR2_X2 U532 ( .A(G146), .B(G125), .ZN(n506) );
  XNOR2_X2 U533 ( .A(n407), .B(G101), .ZN(n505) );
  XNOR2_X2 U534 ( .A(n408), .B(KEYINPUT64), .ZN(n504) );
  XNOR2_X2 U535 ( .A(n409), .B(KEYINPUT45), .ZN(n748) );
  XNOR2_X1 U536 ( .A(n410), .B(n425), .ZN(n497) );
  XNOR2_X2 U537 ( .A(n754), .B(n455), .ZN(n410) );
  INV_X1 U538 ( .A(n573), .ZN(n412) );
  NAND2_X1 U539 ( .A1(n414), .A2(n620), .ZN(n621) );
  XNOR2_X1 U540 ( .A(n416), .B(KEYINPUT122), .ZN(n668) );
  INV_X1 U541 ( .A(n580), .ZN(n418) );
  NAND2_X1 U542 ( .A1(n421), .A2(n712), .ZN(n420) );
  XNOR2_X1 U543 ( .A(n579), .B(KEYINPUT104), .ZN(n421) );
  NAND2_X1 U544 ( .A1(n497), .A2(n496), .ZN(n499) );
  XNOR2_X1 U545 ( .A(n426), .B(n495), .ZN(n425) );
  XNOR2_X1 U546 ( .A(n494), .B(KEYINPUT89), .ZN(n426) );
  XNOR2_X2 U547 ( .A(n530), .B(n434), .ZN(n754) );
  AND2_X2 U548 ( .A1(n656), .A2(n630), .ZN(n509) );
  XNOR2_X2 U549 ( .A(n429), .B(G119), .ZN(n500) );
  NAND2_X1 U550 ( .A1(n433), .A2(n603), .ZN(n432) );
  NAND2_X1 U551 ( .A1(n445), .A2(n374), .ZN(n645) );
  XNOR2_X1 U552 ( .A(n599), .B(KEYINPUT102), .ZN(n445) );
  INV_X1 U553 ( .A(n497), .ZN(n676) );
  NOR2_X1 U554 ( .A1(n585), .A2(n439), .ZN(n438) );
  NAND2_X1 U555 ( .A1(n440), .A2(n449), .ZN(n446) );
  AND2_X1 U556 ( .A1(n440), .A2(KEYINPUT2), .ZN(n737) );
  XNOR2_X1 U557 ( .A(n451), .B(n450), .ZN(G60) );
  NAND2_X1 U558 ( .A1(n452), .A2(n670), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n635), .B(n634), .ZN(n452) );
  XNOR2_X2 U560 ( .A(n509), .B(n508), .ZN(n547) );
  OR2_X2 U561 ( .A1(n709), .A2(n708), .ZN(n711) );
  BUF_X1 U562 ( .A(n667), .Z(n672) );
  XOR2_X2 U563 ( .A(G110), .B(G104), .Z(n502) );
  NOR2_X2 U564 ( .A1(n547), .A2(n577), .ZN(n548) );
  XNOR2_X2 U565 ( .A(n548), .B(KEYINPUT83), .ZN(n554) );
  XNOR2_X2 U566 ( .A(n499), .B(n498), .ZN(n573) );
  INV_X1 U567 ( .A(KEYINPUT79), .ZN(n537) );
  NAND2_X1 U568 ( .A1(n616), .A2(n615), .ZN(n600) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U570 ( .A(n539), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n523), .B(n632), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n505), .B(G146), .ZN(n455) );
  XNOR2_X1 U573 ( .A(n457), .B(n456), .ZN(n462) );
  NAND2_X1 U574 ( .A1(n511), .A2(G210), .ZN(n459) );
  XNOR2_X1 U575 ( .A(n500), .B(n460), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X2 U577 ( .A(n464), .B(G472), .ZN(n543) );
  NAND2_X1 U578 ( .A1(G214), .A2(n507), .ZN(n698) );
  NAND2_X1 U579 ( .A1(n543), .A2(n698), .ZN(n465) );
  XNOR2_X1 U580 ( .A(n466), .B(KEYINPUT87), .ZN(n467) );
  XOR2_X1 U581 ( .A(KEYINPUT14), .B(n467), .Z(n469) );
  NAND2_X1 U582 ( .A1(n469), .A2(G952), .ZN(n468) );
  XOR2_X1 U583 ( .A(KEYINPUT88), .B(n468), .Z(n728) );
  NAND2_X1 U584 ( .A1(n758), .A2(n728), .ZN(n589) );
  NAND2_X1 U585 ( .A1(G902), .A2(n469), .ZN(n587) );
  NOR2_X1 U586 ( .A1(G900), .A2(n587), .ZN(n470) );
  NAND2_X1 U587 ( .A1(G953), .A2(n470), .ZN(n471) );
  NAND2_X1 U588 ( .A1(n589), .A2(n471), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n526), .A2(G221), .ZN(n476) );
  XNOR2_X1 U590 ( .A(n476), .B(n475), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n482) );
  INV_X1 U592 ( .A(G140), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n506), .B(KEYINPUT10), .ZN(n521) );
  NAND2_X1 U596 ( .A1(n630), .A2(G234), .ZN(n486) );
  XNOR2_X1 U597 ( .A(n486), .B(KEYINPUT20), .ZN(n490) );
  NAND2_X1 U598 ( .A1(n490), .A2(G217), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n487), .B(KEYINPUT25), .ZN(n488) );
  NAND2_X1 U600 ( .A1(n490), .A2(G221), .ZN(n492) );
  INV_X1 U601 ( .A(KEYINPUT21), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n594) );
  INV_X1 U603 ( .A(n594), .ZN(n708) );
  NAND2_X1 U604 ( .A1(n758), .A2(G227), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n493), .B(n502), .ZN(n494) );
  XOR2_X1 U606 ( .A(G107), .B(n522), .Z(n495) );
  XNOR2_X1 U607 ( .A(KEYINPUT71), .B(G469), .ZN(n498) );
  XOR2_X2 U608 ( .A(G113), .B(G122), .Z(n510) );
  XOR2_X1 U609 ( .A(n502), .B(n510), .Z(n503) );
  AND2_X1 U610 ( .A1(n507), .A2(G210), .ZN(n508) );
  XOR2_X1 U611 ( .A(n510), .B(KEYINPUT96), .Z(n513) );
  NAND2_X1 U612 ( .A1(G214), .A2(n511), .ZN(n512) );
  XNOR2_X1 U613 ( .A(n513), .B(n512), .ZN(n520) );
  XNOR2_X1 U614 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U615 ( .A(n522), .B(n521), .Z(n753) );
  XNOR2_X1 U616 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n523) );
  INV_X1 U617 ( .A(G475), .ZN(n632) );
  INV_X1 U618 ( .A(n538), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n529), .B(n528), .ZN(n532) );
  INV_X1 U620 ( .A(n530), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U622 ( .A(n534), .B(n533), .ZN(n662) );
  NAND2_X1 U623 ( .A1(n662), .A2(n496), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n535), .B(G478), .ZN(n570) );
  INV_X1 U625 ( .A(n570), .ZN(n558) );
  NOR2_X1 U626 ( .A1(n536), .A2(n558), .ZN(n603) );
  XNOR2_X1 U627 ( .A(n646), .B(n537), .ZN(n552) );
  NAND2_X1 U628 ( .A1(n539), .A2(n594), .ZN(n541) );
  INV_X1 U629 ( .A(KEYINPUT70), .ZN(n540) );
  XNOR2_X1 U630 ( .A(n541), .B(n540), .ZN(n542) );
  AND2_X1 U631 ( .A1(n542), .A2(n709), .ZN(n555) );
  NAND2_X1 U632 ( .A1(n688), .A2(n555), .ZN(n545) );
  BUF_X2 U633 ( .A(n543), .Z(n718) );
  XOR2_X1 U634 ( .A(KEYINPUT6), .B(KEYINPUT101), .Z(n544) );
  NOR2_X1 U635 ( .A1(n545), .A2(n611), .ZN(n546) );
  XNOR2_X1 U636 ( .A(n546), .B(KEYINPUT103), .ZN(n578) );
  INV_X1 U637 ( .A(n698), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n549), .B(KEYINPUT36), .ZN(n551) );
  XOR2_X1 U639 ( .A(KEYINPUT85), .B(n402), .Z(n607) );
  XNOR2_X1 U640 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n718), .A2(n555), .ZN(n557) );
  XNOR2_X1 U642 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n556) );
  OR2_X1 U643 ( .A1(n538), .A2(n558), .ZN(n583) );
  INV_X1 U644 ( .A(n583), .ZN(n690) );
  NOR2_X1 U645 ( .A1(n690), .A2(n688), .ZN(n703) );
  NAND2_X1 U646 ( .A1(n703), .A2(KEYINPUT78), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n639), .A2(n559), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n560), .A2(KEYINPUT47), .ZN(n564) );
  NAND2_X1 U649 ( .A1(n703), .A2(KEYINPUT47), .ZN(n562) );
  INV_X1 U650 ( .A(KEYINPUT78), .ZN(n561) );
  NAND2_X1 U651 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U652 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U653 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n567) );
  NOR2_X1 U654 ( .A1(n703), .A2(n567), .ZN(n568) );
  AND2_X1 U655 ( .A1(n639), .A2(n568), .ZN(n569) );
  INV_X1 U656 ( .A(n576), .ZN(n699) );
  NAND2_X1 U657 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U658 ( .A1(n538), .A2(n570), .ZN(n593) );
  INV_X1 U659 ( .A(n593), .ZN(n701) );
  XOR2_X1 U660 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n571) );
  OR2_X1 U661 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n579) );
  BUF_X1 U663 ( .A(n581), .Z(n582) );
  INV_X1 U664 ( .A(n582), .ZN(n584) );
  NOR2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n641) );
  OR2_X1 U666 ( .A1(n696), .A2(n641), .ZN(n585) );
  NOR2_X1 U667 ( .A1(G898), .A2(n758), .ZN(n743) );
  INV_X1 U668 ( .A(n587), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n743), .A2(n588), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U672 ( .A(n718), .ZN(n620) );
  INV_X1 U673 ( .A(n711), .ZN(n616) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT33), .ZN(n697) );
  INV_X1 U675 ( .A(n611), .ZN(n605) );
  INV_X1 U676 ( .A(n709), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  INV_X1 U679 ( .A(KEYINPUT32), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n402), .A2(n709), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n377), .A2(n613), .ZN(n681) );
  INV_X1 U683 ( .A(n402), .ZN(n712) );
  NAND2_X1 U684 ( .A1(n718), .A2(n616), .ZN(n617) );
  NOR2_X1 U685 ( .A1(n712), .A2(n617), .ZN(n721) );
  NAND2_X1 U686 ( .A1(n721), .A2(n618), .ZN(n619) );
  XNOR2_X1 U687 ( .A(KEYINPUT31), .B(n619), .ZN(n691) );
  NOR2_X1 U688 ( .A1(n376), .A2(n621), .ZN(n684) );
  NOR2_X1 U689 ( .A1(n691), .A2(n684), .ZN(n622) );
  NOR2_X1 U690 ( .A1(n703), .A2(n622), .ZN(n623) );
  NOR2_X1 U691 ( .A1(n681), .A2(n623), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n627), .A2(n748), .ZN(n625) );
  XOR2_X1 U693 ( .A(KEYINPUT80), .B(n630), .Z(n626) );
  INV_X1 U694 ( .A(n630), .ZN(n631) );
  NOR2_X1 U695 ( .A1(n647), .A2(n632), .ZN(n635) );
  XOR2_X1 U696 ( .A(n633), .B(KEYINPUT59), .Z(n634) );
  INV_X1 U697 ( .A(G952), .ZN(n636) );
  NAND2_X1 U698 ( .A1(n636), .A2(G953), .ZN(n670) );
  NAND2_X1 U699 ( .A1(n639), .A2(n690), .ZN(n638) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .Z(n637) );
  XNOR2_X1 U701 ( .A(n638), .B(n637), .ZN(G30) );
  NAND2_X1 U702 ( .A1(n639), .A2(n688), .ZN(n640) );
  XNOR2_X1 U703 ( .A(n640), .B(G146), .ZN(G48) );
  XOR2_X1 U704 ( .A(G134), .B(KEYINPUT111), .Z(n642) );
  XOR2_X1 U705 ( .A(n642), .B(n641), .Z(G36) );
  XOR2_X1 U706 ( .A(G131), .B(n643), .Z(G33) );
  XOR2_X1 U707 ( .A(G110), .B(KEYINPUT109), .Z(n644) );
  XNOR2_X1 U708 ( .A(n645), .B(n644), .ZN(G12) );
  XNOR2_X1 U709 ( .A(n646), .B(G143), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n667), .A2(G472), .ZN(n650) );
  XOR2_X1 U711 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  XNOR2_X1 U712 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U713 ( .A1(n651), .A2(n670), .ZN(n652) );
  XNOR2_X1 U714 ( .A(n652), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n667), .A2(G210), .ZN(n658) );
  XNOR2_X1 U716 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n654) );
  XNOR2_X1 U717 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n653) );
  XNOR2_X1 U718 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U719 ( .A(n381), .B(n655), .ZN(n657) );
  XNOR2_X1 U720 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U721 ( .A1(n659), .A2(n670), .ZN(n661) );
  XOR2_X1 U722 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n660) );
  XNOR2_X1 U723 ( .A(n661), .B(n660), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n667), .A2(G478), .ZN(n664) );
  XNOR2_X1 U725 ( .A(n662), .B(KEYINPUT120), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U727 ( .A1(n665), .A2(n670), .ZN(n666) );
  XNOR2_X1 U728 ( .A(n666), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U729 ( .A1(n672), .A2(G217), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n669), .B(n668), .ZN(n671) );
  INV_X1 U731 ( .A(n670), .ZN(n679) );
  NOR2_X1 U732 ( .A1(n671), .A2(n679), .ZN(G66) );
  NAND2_X1 U733 ( .A1(n672), .A2(G469), .ZN(n678) );
  XNOR2_X1 U734 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n674) );
  XNOR2_X1 U735 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n673) );
  XNOR2_X1 U736 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U737 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U738 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(G54) );
  XOR2_X1 U740 ( .A(G101), .B(n681), .Z(G3) );
  NAND2_X1 U741 ( .A1(n684), .A2(n688), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n682), .B(KEYINPUT108), .ZN(n683) );
  XNOR2_X1 U743 ( .A(G104), .B(n683), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U745 ( .A1(n684), .A2(n690), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U747 ( .A(G107), .B(n687), .ZN(G9) );
  NAND2_X1 U748 ( .A1(n691), .A2(n688), .ZN(n689) );
  XNOR2_X1 U749 ( .A(n689), .B(G113), .ZN(G15) );
  NAND2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n692), .B(G116), .ZN(G18) );
  XOR2_X1 U752 ( .A(KEYINPUT110), .B(KEYINPUT37), .Z(n693) );
  XNOR2_X1 U753 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U754 ( .A(G125), .B(n695), .ZN(G27) );
  XOR2_X1 U755 ( .A(G140), .B(n696), .Z(G42) );
  XNOR2_X1 U756 ( .A(KEYINPUT115), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT114), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n731), .A2(n707), .ZN(n725) );
  NAND2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U764 ( .A(KEYINPUT49), .B(n710), .Z(n716) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n713), .B(KEYINPUT50), .ZN(n714) );
  XNOR2_X1 U767 ( .A(KEYINPUT112), .B(n714), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U770 ( .A(KEYINPUT113), .B(n719), .Z(n720) );
  NOR2_X1 U771 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U772 ( .A(KEYINPUT51), .B(n722), .Z(n723) );
  NOR2_X1 U773 ( .A1(n730), .A2(n723), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n729) );
  AND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(n733) );
  NOR2_X1 U777 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U778 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U779 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U780 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U781 ( .A(KEYINPUT116), .B(n738), .Z(n739) );
  NOR2_X1 U782 ( .A1(G953), .A2(n739), .ZN(n740) );
  XNOR2_X1 U783 ( .A(KEYINPUT53), .B(n740), .ZN(G75) );
  XOR2_X1 U784 ( .A(n741), .B(G101), .Z(n742) );
  NOR2_X1 U785 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U786 ( .A(KEYINPUT124), .B(n744), .Z(n752) );
  XOR2_X1 U787 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n746) );
  NAND2_X1 U788 ( .A1(G224), .A2(G953), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n746), .B(n745), .ZN(n747) );
  NAND2_X1 U790 ( .A1(n747), .A2(G898), .ZN(n750) );
  NAND2_X1 U791 ( .A1(n379), .A2(n758), .ZN(n749) );
  NAND2_X1 U792 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U793 ( .A(n752), .B(n751), .Z(G69) );
  XNOR2_X1 U794 ( .A(n753), .B(KEYINPUT125), .ZN(n755) );
  XNOR2_X1 U795 ( .A(n754), .B(n755), .ZN(n760) );
  INV_X1 U796 ( .A(n760), .ZN(n756) );
  XNOR2_X1 U797 ( .A(n756), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U798 ( .A(n628), .B(n757), .ZN(n759) );
  NAND2_X1 U799 ( .A1(n759), .A2(n758), .ZN(n764) );
  XNOR2_X1 U800 ( .A(G227), .B(n760), .ZN(n761) );
  NAND2_X1 U801 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U802 ( .A1(n762), .A2(G953), .ZN(n763) );
  NAND2_X1 U803 ( .A1(n764), .A2(n763), .ZN(G72) );
  XNOR2_X1 U804 ( .A(n765), .B(n528), .ZN(n766) );
  XNOR2_X1 U805 ( .A(n766), .B(KEYINPUT127), .ZN(G24) );
  BUF_X1 U806 ( .A(n767), .Z(n768) );
  XNOR2_X1 U807 ( .A(G119), .B(n768), .ZN(G21) );
  XOR2_X1 U808 ( .A(n769), .B(G137), .Z(G39) );
endmodule

