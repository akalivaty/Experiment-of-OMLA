//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n450), .B(new_n451), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  INV_X1    g054(.A(G138), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n463), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT4), .B1(new_n481), .B2(KEYINPUT67), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n464), .A2(G138), .A3(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .A3(new_n484), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n474), .B2(G126), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT69), .Z(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n503), .A2(new_n515), .ZN(G166));
  NOR2_X1   g091(.A1(new_n510), .A2(new_n509), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n504), .B2(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n513), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n523), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n521), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n498), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n535), .B2(new_n534), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n539));
  INV_X1    g114(.A(new_n513), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G90), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n541), .B1(G52), .B2(new_n525), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n507), .A2(new_n545), .B1(new_n513), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n521), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(KEYINPUT74), .A3(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n547), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n525), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT75), .B(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n517), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G651), .A2(new_n565), .B1(new_n540), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  INV_X1    g144(.A(G49), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n507), .A2(new_n570), .B1(new_n513), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n522), .A2(G74), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(G651), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n498), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n507), .A2(new_n578), .B1(new_n513), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n521), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n540), .A2(G85), .B1(G47), .B2(new_n525), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n506), .A2(new_n501), .A3(KEYINPUT10), .A4(G92), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(G66), .B1(new_n510), .B2(new_n509), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n598), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT77), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n598), .A2(new_n602), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n598), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n608), .A2(KEYINPUT78), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n592), .B1(G868), .B2(new_n611), .ZN(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n611), .B2(new_n618), .ZN(new_n621));
  AOI211_X1 g196(.A(KEYINPUT80), .B(G559), .C1(new_n605), .C2(new_n610), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n621), .A2(new_n622), .A3(new_n614), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n614), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n464), .A2(new_n469), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n468), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n474), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n466), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G6), .A2(G16), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n581), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n574), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n690), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n689), .A2(new_n695), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT85), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT85), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT86), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(new_n702), .B2(new_n703), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n589), .A2(new_n590), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n690), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n690), .B2(G24), .ZN(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n468), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n474), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(new_n714), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT83), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n711), .A2(new_n712), .ZN(new_n726));
  NOR4_X1   g301(.A1(new_n708), .A2(new_n713), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n707), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n707), .B2(new_n727), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n690), .A2(G20), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT23), .Z(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1956), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G160), .A2(G29), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NOR2_X1   g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n714), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT93), .ZN(new_n742));
  AOI21_X1  g317(.A(G2084), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT96), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G28), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n714), .B1(new_n746), .B2(G28), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n745), .B1(new_n747), .B2(new_n748), .C1(new_n636), .C2(new_n714), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n714), .A2(G32), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  INV_X1    g330(.A(new_n474), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n714), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n738), .A2(G2084), .A3(new_n742), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n714), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n468), .A2(G140), .ZN(new_n767));
  INV_X1    g342(.A(G128), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n756), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G116), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT89), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(new_n714), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT90), .B(G2067), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n750), .A2(new_n763), .A3(new_n764), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n714), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n714), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT29), .Z(new_n782));
  AOI211_X1 g357(.A(new_n737), .B(new_n778), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G168), .A2(G16), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(KEYINPUT95), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT95), .B2(new_n784), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1966), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2072), .ZN(new_n790));
  OR2_X1    g365(.A1(G29), .A2(G33), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n468), .A2(G139), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT91), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT91), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(G115), .A2(G2104), .ZN(new_n797));
  INV_X1    g372(.A(G127), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n463), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(KEYINPUT92), .B1(new_n799), .B2(G2105), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n799), .A2(KEYINPUT92), .A3(G2105), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n795), .A2(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n791), .B1(new_n802), .B2(new_n714), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n782), .A2(new_n779), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n790), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n555), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G16), .B2(G19), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT88), .B(G1341), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G27), .A2(G29), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G164), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2078), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n807), .A2(new_n808), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n805), .A2(new_n809), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G5), .A2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G301), .B2(new_n690), .ZN(new_n817));
  INV_X1    g392(.A(G1961), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NOR2_X1   g395(.A1(G4), .A2(G16), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n611), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n789), .A2(new_n814), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n731), .A2(new_n732), .A3(new_n827), .ZN(G311));
  NOR2_X1   g403(.A1(new_n732), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n730), .ZN(G150));
  NAND3_X1  g405(.A1(new_n519), .A2(new_n520), .A3(G67), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G651), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n540), .A2(G93), .B1(G55), .B2(new_n525), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n834), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n611), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n840), .A2(new_n555), .A3(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n553), .A2(new_n554), .ZN(new_n846));
  INV_X1    g421(.A(new_n547), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n836), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(KEYINPUT99), .C1(new_n840), .C2(new_n555), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n844), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT100), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(KEYINPUT100), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n842), .B1(new_n855), .B2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n471), .B(new_n636), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n478), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n496), .A2(KEYINPUT101), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n487), .A2(new_n491), .A3(new_n862), .A4(new_n495), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n468), .A2(G142), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n474), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n466), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n627), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n802), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n759), .ZN(new_n874));
  INV_X1    g449(.A(new_n759), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n802), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n720), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n720), .A3(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(new_n871), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n865), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n881), .B2(new_n877), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n879), .A3(new_n871), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n864), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n887), .A3(new_n774), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n774), .B1(new_n884), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n860), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(KEYINPUT104), .A3(new_n859), .A4(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(G290), .A2(G288), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n709), .A2(new_n574), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  XOR2_X1   g477(.A(G166), .B(new_n581), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n900), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n906), .A2(KEYINPUT106), .A3(new_n903), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n904), .ZN(new_n909));
  INV_X1    g484(.A(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  INV_X1    g487(.A(new_n907), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n621), .B2(new_n622), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n603), .A2(new_n604), .A3(new_n593), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT78), .B1(new_n608), .B2(new_n609), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n618), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT80), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n611), .A2(new_n620), .A3(new_n618), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT105), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n917), .A2(new_n923), .A3(new_n850), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n850), .B1(new_n917), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g500(.A(G299), .B(new_n606), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n850), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n621), .A2(new_n622), .A3(new_n916), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n921), .B2(new_n922), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n917), .A2(new_n923), .A3(new_n850), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT107), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n926), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n924), .B2(new_n925), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n934), .A3(new_n927), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n915), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n915), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n840), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(G868), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(G295));
  AND2_X1   g523(.A1(new_n908), .A2(new_n914), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n938), .A2(new_n940), .A3(new_n939), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n915), .A2(new_n941), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n614), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n954), .A2(KEYINPUT108), .A3(new_n946), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n944), .B2(new_n947), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(G331));
  AND3_X1   g533(.A1(new_n845), .A2(new_n849), .A3(G286), .ZN(new_n959));
  AOI21_X1  g534(.A(G286), .B1(new_n845), .B2(new_n849), .ZN(new_n960));
  OAI21_X1  g535(.A(G301), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n850), .A2(G168), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n845), .A2(new_n849), .A3(G286), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(G171), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n961), .A2(new_n964), .A3(new_n927), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n926), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n965), .A2(new_n966), .B1(new_n907), .B2(new_n905), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n905), .A2(new_n907), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n964), .A3(new_n927), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n961), .A2(new_n964), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n926), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n967), .A2(new_n971), .A3(new_n976), .A4(new_n895), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n967), .A2(new_n971), .A3(new_n895), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n967), .A2(new_n971), .A3(new_n976), .A4(new_n972), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n978), .A2(new_n982), .ZN(G397));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n861), .A2(new_n984), .A3(new_n863), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n467), .A2(G40), .A3(new_n470), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n774), .B(G2067), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n759), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n720), .A2(new_n724), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n720), .A2(new_n724), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n998), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n709), .A2(new_n712), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n989), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n997), .A2(new_n998), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n990), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n990), .B1(new_n875), .B2(new_n992), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n990), .B2(new_n993), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n989), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1009), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n988), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n496), .A2(new_n984), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n986), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n496), .A2(new_n1026), .A3(KEYINPUT45), .A4(new_n984), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1023), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n496), .A2(new_n1034), .A3(new_n984), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT110), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n496), .A2(new_n1037), .A3(new_n1034), .A4(new_n984), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT116), .B(G2084), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1032), .A2(G168), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(KEYINPUT120), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(G8), .A3(G286), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1042), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT62), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n984), .A4(new_n863), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1025), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n698), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1033), .A2(new_n1036), .A3(new_n779), .A4(new_n1038), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G166), .A2(new_n1043), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(KEYINPUT111), .B2(KEYINPUT55), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n496), .A2(new_n984), .A3(new_n988), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n574), .A2(G1976), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n574), .B2(G1976), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1061), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT113), .B(G1981), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n581), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n688), .B2(new_n581), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1060), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1033), .A2(new_n779), .A3(new_n1035), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1971), .B1(new_n1025), .B2(new_n1051), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1059), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1052), .B2(G2078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT122), .B(G1961), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1087), .A2(G2078), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1025), .A2(new_n1029), .A3(new_n1027), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1080), .A2(new_n1086), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1047), .A4(new_n1045), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1050), .A2(new_n1096), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1043), .B(G286), .C1(new_n1032), .C2(new_n1040), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(new_n1085), .A3(new_n1060), .A4(new_n1079), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND4_X1   g680(.A1(KEYINPUT63), .A2(new_n1046), .A3(G8), .A4(G168), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1078), .B1(new_n1059), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1084), .B1(new_n1107), .B2(KEYINPUT117), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1106), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1060), .A2(new_n1078), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT114), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1074), .B1(new_n1115), .B2(new_n1076), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1072), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1101), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(G299), .B(KEYINPUT57), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n736), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT56), .B(G2072), .Z(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1025), .A2(new_n1051), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1119), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1119), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1120), .B2(new_n736), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n1124), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT119), .B1(new_n1132), .B2(KEYINPUT61), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1125), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1131), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1061), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1089), .A2(new_n823), .B1(new_n1010), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n603), .A2(new_n604), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1128), .A2(KEYINPUT61), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n1125), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT58), .B(G1341), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1052), .A2(G1996), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n555), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1148), .B2(new_n555), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1143), .B1(new_n1142), .B2(KEYINPUT60), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1133), .A2(new_n1140), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1134), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1051), .A2(new_n1092), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n988), .B(KEYINPUT124), .Z(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n985), .B2(new_n986), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1091), .B(KEYINPUT123), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(G301), .A4(new_n1088), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1160), .B1(new_n1168), .B2(new_n1095), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT54), .B1(new_n1094), .B2(G171), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1166), .A2(new_n1167), .A3(new_n1088), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(G171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1085), .B(new_n1108), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1118), .B1(new_n1159), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n989), .B1(new_n1006), .B2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1002), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1022), .B1(new_n1175), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g754(.A1(new_n974), .A2(new_n977), .ZN(new_n1181));
  NOR4_X1   g755(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n896), .A3(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


