

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591;

  NAND2_X1 U321 ( .A1(n578), .A2(n561), .ZN(n359) );
  INV_X1 U322 ( .A(n570), .ZN(n481) );
  NOR2_X2 U323 ( .A1(n527), .A2(n424), .ZN(n577) );
  XOR2_X1 U324 ( .A(n331), .B(n330), .Z(n578) );
  XOR2_X1 U325 ( .A(n428), .B(n368), .Z(n289) );
  INV_X1 U326 ( .A(n498), .ZN(n394) );
  AND2_X1 U327 ( .A1(n396), .A2(n395), .ZN(n398) );
  XNOR2_X1 U328 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  INV_X1 U329 ( .A(KEYINPUT48), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n337), .B(n336), .ZN(n415) );
  XNOR2_X1 U331 ( .A(n406), .B(n405), .ZN(n539) );
  XNOR2_X1 U332 ( .A(n358), .B(n357), .ZN(n582) );
  XOR2_X1 U333 ( .A(n377), .B(n376), .Z(n570) );
  XOR2_X1 U334 ( .A(n312), .B(n311), .Z(n527) );
  XNOR2_X1 U335 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U336 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n442) );
  XOR2_X1 U338 ( .A(KEYINPUT3), .B(KEYINPUT88), .Z(n291) );
  XNOR2_X1 U339 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n435) );
  XOR2_X1 U341 ( .A(n435), .B(KEYINPUT91), .Z(n293) );
  NAND2_X1 U342 ( .A1(G225GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n312) );
  XOR2_X1 U344 ( .A(G57GAT), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U345 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n297) );
  XNOR2_X1 U348 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(n299), .B(n298), .Z(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U352 ( .A(KEYINPUT83), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(G113GAT), .B(n302), .Z(n453) );
  XOR2_X1 U355 ( .A(G85GAT), .B(G155GAT), .Z(n304) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G148GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT78), .Z(n365) );
  XOR2_X1 U359 ( .A(n305), .B(n365), .Z(n307) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G162GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n453), .B(n308), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U364 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n314) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(KEYINPUT67), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n331) );
  XOR2_X1 U367 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n373) );
  XNOR2_X1 U370 ( .A(G15GAT), .B(G1GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n317), .B(G8GAT), .ZN(n382) );
  XNOR2_X1 U372 ( .A(n373), .B(n382), .ZN(n321) );
  XNOR2_X1 U373 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(KEYINPUT29), .ZN(n319) );
  XOR2_X1 U375 ( .A(n319), .B(KEYINPUT30), .Z(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n327) );
  XOR2_X1 U377 ( .A(G113GAT), .B(G22GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G141GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U380 ( .A(G50GAT), .B(G36GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  INV_X1 U385 ( .A(G92GAT), .ZN(n332) );
  NAND2_X1 U386 ( .A1(G64GAT), .A2(n332), .ZN(n335) );
  INV_X1 U387 ( .A(G64GAT), .ZN(n333) );
  NAND2_X1 U388 ( .A1(n333), .A2(G92GAT), .ZN(n334) );
  NAND2_X1 U389 ( .A1(n335), .A2(n334), .ZN(n337) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  INV_X1 U391 ( .A(n446), .ZN(n338) );
  NAND2_X1 U392 ( .A1(n415), .A2(n338), .ZN(n341) );
  INV_X1 U393 ( .A(n415), .ZN(n339) );
  NAND2_X1 U394 ( .A1(n339), .A2(n446), .ZN(n340) );
  NAND2_X1 U395 ( .A1(n341), .A2(n340), .ZN(n343) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n344), .B(KEYINPUT71), .ZN(n348) );
  INV_X1 U399 ( .A(n348), .ZN(n346) );
  XOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT13), .Z(n381) );
  XOR2_X1 U401 ( .A(n381), .B(KEYINPUT70), .Z(n347) );
  INV_X1 U402 ( .A(n347), .ZN(n345) );
  NAND2_X1 U403 ( .A1(n346), .A2(n345), .ZN(n350) );
  NAND2_X1 U404 ( .A1(n348), .A2(n347), .ZN(n349) );
  NAND2_X1 U405 ( .A1(n350), .A2(n349), .ZN(n354) );
  XOR2_X1 U406 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n352) );
  XNOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n351) );
  XOR2_X1 U408 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n358) );
  XNOR2_X1 U410 ( .A(G106GAT), .B(G78GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n355), .B(G148GAT), .ZN(n437) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G85GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n356), .B(KEYINPUT72), .ZN(n368) );
  XNOR2_X1 U414 ( .A(n437), .B(n368), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n582), .B(KEYINPUT41), .ZN(n561) );
  XNOR2_X1 U416 ( .A(n359), .B(KEYINPUT46), .ZN(n396) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT76), .B(KEYINPUT64), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n377) );
  XOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n363) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(G92GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U423 ( .A(n364), .B(KEYINPUT9), .Z(n367) );
  XNOR2_X1 U424 ( .A(G218GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U426 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n289), .B(n369), .ZN(n370) );
  XOR2_X1 U429 ( .A(n371), .B(n370), .Z(n375) );
  XNOR2_X1 U430 ( .A(G36GAT), .B(G190GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n372), .B(KEYINPUT79), .ZN(n417) );
  XNOR2_X1 U432 ( .A(n373), .B(n417), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U434 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n379) );
  XNOR2_X1 U435 ( .A(G183GAT), .B(G64GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n384) );
  XOR2_X1 U438 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XNOR2_X1 U439 ( .A(n382), .B(n427), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n386) );
  NAND2_X1 U442 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U444 ( .A(n388), .B(n387), .Z(n393) );
  XOR2_X1 U445 ( .A(G78GAT), .B(G211GAT), .Z(n390) );
  XNOR2_X1 U446 ( .A(G127GAT), .B(G71GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n391), .B(KEYINPUT12), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n498) );
  NOR2_X1 U450 ( .A1(n570), .A2(n394), .ZN(n395) );
  XNOR2_X1 U451 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n404) );
  XNOR2_X1 U453 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT36), .B(n481), .ZN(n588) );
  NOR2_X1 U455 ( .A1(n588), .A2(n498), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U457 ( .A1(n401), .A2(n578), .ZN(n402) );
  NAND2_X1 U458 ( .A1(n582), .A2(n402), .ZN(n403) );
  NAND2_X1 U459 ( .A1(n404), .A2(n403), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n408) );
  XNOR2_X1 U461 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U463 ( .A(G169GAT), .B(n409), .Z(n452) );
  XOR2_X1 U464 ( .A(KEYINPUT87), .B(G218GAT), .Z(n411) );
  XNOR2_X1 U465 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U467 ( .A(G197GAT), .B(n412), .Z(n438) );
  XNOR2_X1 U468 ( .A(n452), .B(n438), .ZN(n421) );
  XOR2_X1 U469 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n414) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U472 ( .A(n416), .B(n415), .Z(n419) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n529) );
  XNOR2_X1 U476 ( .A(n529), .B(KEYINPUT121), .ZN(n422) );
  NOR2_X1 U477 ( .A1(n539), .A2(n422), .ZN(n423) );
  XOR2_X1 U478 ( .A(KEYINPUT54), .B(n423), .Z(n424) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U480 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n477) );
  NAND2_X1 U491 ( .A1(n577), .A2(n477), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n458) );
  XOR2_X1 U493 ( .A(G176GAT), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(G134GAT), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U496 ( .A(n445), .B(G190GAT), .Z(n448) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n457) );
  XOR2_X1 U499 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n450) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U502 ( .A(n451), .B(KEYINPUT20), .Z(n455) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U505 ( .A(n457), .B(n456), .Z(n467) );
  NOR2_X2 U506 ( .A1(n458), .A2(n467), .ZN(n460) );
  INV_X1 U507 ( .A(KEYINPUT123), .ZN(n459) );
  XNOR2_X2 U508 ( .A(n460), .B(n459), .ZN(n571) );
  NAND2_X1 U509 ( .A1(n571), .A2(n578), .ZN(n462) );
  XNOR2_X1 U510 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n462), .B(n461), .ZN(G1348GAT) );
  NAND2_X1 U512 ( .A1(n571), .A2(n561), .ZN(n465) );
  XOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n487) );
  NAND2_X1 U515 ( .A1(n582), .A2(n578), .ZN(n466) );
  XNOR2_X1 U516 ( .A(n466), .B(KEYINPUT74), .ZN(n502) );
  INV_X1 U517 ( .A(n467), .ZN(n540) );
  NAND2_X1 U518 ( .A1(n529), .A2(n540), .ZN(n468) );
  NAND2_X1 U519 ( .A1(n468), .A2(n477), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT96), .B(n469), .Z(n470) );
  XNOR2_X1 U521 ( .A(n470), .B(KEYINPUT25), .ZN(n473) );
  NOR2_X1 U522 ( .A1(n540), .A2(n477), .ZN(n471) );
  XNOR2_X1 U523 ( .A(n471), .B(KEYINPUT26), .ZN(n576) );
  XNOR2_X1 U524 ( .A(n529), .B(KEYINPUT27), .ZN(n476) );
  NAND2_X1 U525 ( .A1(n576), .A2(n476), .ZN(n472) );
  NAND2_X1 U526 ( .A1(n473), .A2(n472), .ZN(n475) );
  INV_X1 U527 ( .A(n527), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n527), .A2(n476), .ZN(n538) );
  NOR2_X1 U530 ( .A1(n540), .A2(n538), .ZN(n478) );
  XNOR2_X1 U531 ( .A(n477), .B(KEYINPUT28), .ZN(n543) );
  NAND2_X1 U532 ( .A1(n478), .A2(n543), .ZN(n479) );
  NAND2_X1 U533 ( .A1(n480), .A2(n479), .ZN(n497) );
  XOR2_X1 U534 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n483) );
  NAND2_X1 U535 ( .A1(n394), .A2(n481), .ZN(n482) );
  XNOR2_X1 U536 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U537 ( .A1(n497), .A2(n484), .ZN(n485) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(n485), .Z(n515) );
  NOR2_X1 U539 ( .A1(n502), .A2(n515), .ZN(n494) );
  NAND2_X1 U540 ( .A1(n494), .A2(n527), .ZN(n486) );
  XNOR2_X1 U541 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  XOR2_X1 U543 ( .A(G8GAT), .B(KEYINPUT99), .Z(n490) );
  NAND2_X1 U544 ( .A1(n494), .A2(n529), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U547 ( .A1(n494), .A2(n540), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  XOR2_X1 U550 ( .A(G22GAT), .B(KEYINPUT101), .Z(n496) );
  INV_X1 U551 ( .A(n543), .ZN(n533) );
  NAND2_X1 U552 ( .A1(n494), .A2(n533), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n496), .B(n495), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n498), .A2(n497), .ZN(n499) );
  NOR2_X1 U555 ( .A1(n588), .A2(n499), .ZN(n500) );
  XOR2_X1 U556 ( .A(KEYINPUT37), .B(n500), .Z(n501) );
  XNOR2_X1 U557 ( .A(KEYINPUT103), .B(n501), .ZN(n526) );
  NOR2_X1 U558 ( .A1(n526), .A2(n502), .ZN(n503) );
  XNOR2_X1 U559 ( .A(n503), .B(KEYINPUT38), .ZN(n512) );
  NAND2_X1 U560 ( .A1(n512), .A2(n527), .ZN(n507) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n505) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U564 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  XOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U566 ( .A1(n529), .A2(n512), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n512), .A2(n540), .ZN(n510) );
  XNOR2_X1 U569 ( .A(n510), .B(KEYINPUT40), .ZN(n511) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n533), .A2(n512), .ZN(n513) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n513), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n517) );
  INV_X1 U574 ( .A(n578), .ZN(n514) );
  NAND2_X1 U575 ( .A1(n514), .A2(n561), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n515), .A2(n525), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n527), .A2(n521), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n521), .A2(n529), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n518), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n540), .A2(n521), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U585 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n527), .A2(n534), .ZN(n528) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(KEYINPUT108), .ZN(n531) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n540), .A2(n534), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n536) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n558) );
  NAND2_X1 U601 ( .A1(n558), .A2(n540), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT112), .B(n541), .Z(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT113), .ZN(n554) );
  NAND2_X1 U605 ( .A1(n578), .A2(n554), .ZN(n545) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U608 ( .A1(n554), .A2(n561), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT114), .Z(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n553) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n551) );
  NAND2_X1 U614 ( .A1(n554), .A2(n394), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U618 ( .A1(n554), .A2(n570), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT119), .ZN(n560) );
  AND2_X1 U622 ( .A1(n558), .A2(n576), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n567), .A2(n578), .ZN(n559) );
  XOR2_X1 U624 ( .A(n560), .B(n559), .Z(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n563) );
  NAND2_X1 U627 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n394), .A2(n567), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n570), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n394), .A2(n571), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n587) );
  INV_X1 U642 ( .A(n587), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n585), .A2(n578), .ZN(n581) );
  XOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .Z(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT59), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  OR2_X1 U648 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n394), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

