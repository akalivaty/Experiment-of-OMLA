//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT80), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(G101), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n193), .A3(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT77), .A2(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT77), .A2(G101), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n195), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(G143), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n209), .A2(new_n210), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n214), .A3(G146), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n207), .A4(G128), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n195), .B(KEYINPUT78), .C1(new_n199), .C2(new_n203), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n206), .A2(new_n221), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n193), .A2(G104), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n201), .ZN(new_n229));
  INV_X1    g043(.A(new_n199), .ZN(new_n230));
  INV_X1    g044(.A(new_n203), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G143), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n233), .B2(G146), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n234), .A2(G128), .B1(new_n222), .B2(new_n223), .ZN(new_n235));
  INV_X1    g049(.A(new_n224), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G134), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n245), .A3(new_n243), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n239), .B2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n246), .ZN(new_n252));
  INV_X1    g066(.A(new_n244), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n257));
  AND4_X1   g071(.A1(new_n190), .A2(new_n238), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n237), .B2(new_n226), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n259), .A2(KEYINPUT12), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n190), .B1(new_n259), .B2(new_n257), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n215), .A2(new_n220), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n222), .A2(new_n223), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n263), .A2(new_n267), .B1(new_n268), .B2(new_n265), .ZN(new_n269));
  OAI21_X1  g083(.A(G101), .B1(new_n199), .B2(new_n194), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n270), .A2(KEYINPUT4), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n230), .A2(new_n231), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(KEYINPUT4), .C1(new_n270), .C2(KEYINPUT76), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n269), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n215), .A2(new_n220), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n210), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n224), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n206), .ZN(new_n279));
  INV_X1    g093(.A(new_n225), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT10), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n237), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n275), .A2(new_n281), .A3(new_n283), .A4(new_n255), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n262), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G110), .B(G140), .ZN(new_n286));
  INV_X1    g100(.A(G227), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n289), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n275), .A2(new_n281), .A3(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n256), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n285), .A2(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n189), .B1(new_n294), .B2(G469), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n284), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n289), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n259), .A2(new_n190), .A3(new_n257), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n238), .A2(new_n256), .A3(new_n257), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT80), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n259), .A2(KEYINPUT12), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT81), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n300), .C1(new_n302), .C2(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(new_n291), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n299), .B1(new_n308), .B2(KEYINPUT82), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n305), .A2(new_n310), .A3(new_n307), .A4(new_n291), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n296), .B1(new_n312), .B2(new_n187), .ZN(new_n313));
  INV_X1    g127(.A(G221), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(new_n188), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n320), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n324), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n326));
  INV_X1    g140(.A(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G116), .ZN(new_n328));
  OAI21_X1  g142(.A(G113), .B1(new_n328), .B2(KEYINPUT5), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n321), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n206), .B2(new_n225), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n332), .A3(new_n334), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT83), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n267), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n222), .A2(new_n223), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n276), .A2(new_n341), .B1(new_n342), .B2(new_n264), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(G125), .B2(new_n278), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT84), .B(G224), .Z(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n333), .B(new_n335), .C1(KEYINPUT83), .C2(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n340), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT7), .B1(new_n346), .B2(G953), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n344), .B(new_n353), .C1(G125), .C2(new_n278), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n334), .B(KEYINPUT8), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n330), .A2(new_n204), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n331), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n337), .A2(new_n352), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n188), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G210), .B1(G237), .B2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n350), .A2(new_n359), .A3(new_n361), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT85), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n366));
  NAND2_X1  g180(.A1(KEYINPUT18), .A2(G131), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G214), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(new_n211), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n233), .A2(new_n370), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(KEYINPUT86), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n375));
  INV_X1    g189(.A(new_n367), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n208), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT73), .A2(G125), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(G146), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n373), .A2(G131), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n371), .A2(new_n372), .A3(new_n250), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(KEYINPUT87), .A3(new_n389), .ZN(new_n390));
  OR3_X1    g204(.A1(new_n373), .A2(KEYINPUT87), .A3(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT19), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n383), .A2(KEYINPUT19), .A3(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n208), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT16), .B1(new_n382), .B2(G125), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT88), .A4(new_n208), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n387), .B1(new_n392), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(G113), .B(G122), .Z(new_n408));
  XOR2_X1   g222(.A(KEYINPUT89), .B(G104), .Z(new_n409));
  XOR2_X1   g223(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT17), .B1(new_n390), .B2(new_n391), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n216), .A3(new_n402), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(new_n404), .C1(new_n388), .C2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n387), .B(new_n410), .C1(new_n413), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n366), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT20), .B(new_n421), .C1(new_n412), .C2(new_n417), .ZN(new_n422));
  INV_X1    g236(.A(G475), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n387), .B1(new_n413), .B2(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n411), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n425), .B2(new_n417), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n420), .A2(new_n422), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G217), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n315), .A2(new_n428), .A3(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n233), .A2(G128), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n210), .A2(G143), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G134), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(KEYINPUT13), .A3(new_n431), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(G134), .C1(KEYINPUT13), .C2(new_n430), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(G107), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n438), .A2(KEYINPUT90), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(KEYINPUT90), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n434), .B(new_n436), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n193), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n193), .B1(new_n446), .B2(KEYINPUT14), .ZN(new_n447));
  AOI22_X1  g261(.A1(KEYINPUT91), .A2(new_n442), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n239), .B1(new_n430), .B2(new_n431), .ZN(new_n449));
  OAI221_X1 g263(.A(new_n448), .B1(KEYINPUT91), .B2(new_n442), .C1(new_n433), .C2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n450), .A3(new_n429), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(KEYINPUT93), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G952), .ZN(new_n463));
  AOI211_X1 g277(.A(G953), .B(new_n463), .C1(G234), .C2(G237), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(G898), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT94), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n188), .B(new_n369), .C1(G234), .C2(G237), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n453), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT93), .B(new_n188), .C1(new_n471), .C2(new_n451), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n427), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n350), .A2(new_n359), .A3(new_n477), .A4(new_n361), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n365), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n313), .A2(new_n317), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n324), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n250), .B1(new_n242), .B2(new_n240), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n249), .B2(new_n250), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n278), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n481), .B(new_n484), .C1(new_n255), .C2(new_n343), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n269), .B1(new_n254), .B2(new_n251), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(KEYINPUT67), .A3(new_n481), .A4(new_n484), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n491), .A3(new_n484), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n488), .B2(new_n484), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n324), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n495));
  NAND3_X1  g309(.A1(new_n368), .A2(new_n369), .A3(G210), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT31), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n490), .A2(new_n494), .A3(KEYINPUT31), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n488), .A2(new_n484), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n324), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n487), .A3(new_n489), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT28), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n485), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(G472), .A2(G902), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT69), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT32), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n517), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT32), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n487), .A2(new_n489), .ZN(new_n525));
  INV_X1    g339(.A(new_n493), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n488), .A2(new_n491), .A3(new_n484), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n525), .B1(new_n528), .B2(new_n324), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n524), .B1(new_n529), .B2(new_n499), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n188), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n499), .A2(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT70), .B1(new_n507), .B2(KEYINPUT28), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n532), .B(new_n533), .C1(new_n511), .C2(KEYINPUT70), .ZN(new_n534));
  OAI21_X1  g348(.A(G472), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n514), .A2(new_n536), .A3(KEYINPUT32), .A4(new_n517), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n519), .A2(new_n522), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n327), .A2(G128), .ZN(new_n539));
  AND2_X1   g353(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n210), .A2(G119), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n544), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n545), .A2(KEYINPUT74), .A3(G110), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n545), .B2(G110), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n539), .A2(new_n543), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT24), .B(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n404), .A3(new_n380), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n404), .A2(new_n414), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(G110), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n555), .C1(new_n549), .C2(new_n550), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n556), .A3(new_n560), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n188), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT25), .Z(new_n565));
  AOI21_X1  g379(.A(new_n428), .B1(G234), .B2(new_n188), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G902), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n567), .B(KEYINPUT75), .Z(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n562), .A2(new_n563), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n565), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n480), .A2(new_n538), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n200), .A2(new_n202), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G3));
  INV_X1    g388(.A(new_n317), .ZN(new_n575));
  AOI211_X1 g389(.A(G469), .B(G902), .C1(new_n309), .C2(new_n311), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(new_n296), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n514), .A2(new_n578), .A3(new_n188), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n502), .A2(new_n503), .B1(new_n511), .B2(new_n512), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT95), .B1(new_n580), .B2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n581), .A3(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n520), .ZN(new_n583));
  INV_X1    g397(.A(new_n571), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n476), .ZN(new_n586));
  INV_X1    g400(.A(new_n363), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(KEYINPUT96), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n363), .A2(new_n589), .A3(new_n364), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT33), .B1(new_n471), .B2(new_n451), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n452), .A2(new_n594), .A3(new_n453), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n455), .A2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT97), .B(G478), .Z(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n454), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n597), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n593), .B2(new_n595), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n454), .A2(new_n600), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n420), .A2(new_n422), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n426), .A2(new_n423), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n603), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n592), .A2(KEYINPUT99), .A3(new_n470), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n470), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n591), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n585), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n422), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n609), .B(new_n620), .C1(new_n608), .C2(new_n619), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n462), .A2(new_n473), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR4_X1   g437(.A1(new_n591), .A2(new_n621), .A3(new_n469), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n585), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n565), .A2(new_n566), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n561), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n557), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n569), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n582), .A2(new_n632), .A3(new_n520), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n582), .A2(new_n632), .A3(KEYINPUT101), .A4(new_n520), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n480), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  AND2_X1   g453(.A1(new_n538), .A2(new_n632), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n577), .A2(new_n591), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n468), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n464), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n621), .A2(new_n623), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XNOR2_X1  g463(.A(new_n645), .B(KEYINPUT39), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OR3_X1    g465(.A1(new_n577), .A2(KEYINPUT40), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT40), .B1(new_n577), .B2(new_n651), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n365), .A2(new_n478), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT38), .Z(new_n655));
  NOR2_X1   g469(.A1(new_n529), .A2(new_n512), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n188), .B1(new_n507), .B2(new_n499), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n519), .A2(new_n522), .A3(new_n537), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n427), .A2(new_n622), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n632), .A2(new_n586), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n652), .A2(new_n653), .A3(new_n655), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(new_n233), .Z(G45));
  INV_X1    g478(.A(new_n632), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n610), .A2(new_n645), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n641), .A2(new_n538), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  NAND2_X1  g483(.A1(new_n538), .A2(new_n571), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n291), .B1(new_n262), .B2(new_n306), .ZN(new_n672));
  INV_X1    g486(.A(new_n307), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT82), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n311), .A3(new_n298), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n188), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n187), .A3(new_n188), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n679));
  OR3_X1    g493(.A1(new_n312), .A2(KEYINPUT102), .A3(new_n187), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n317), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n615), .A2(new_n671), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT103), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n671), .A2(new_n615), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND3_X1  g502(.A1(new_n671), .A2(new_n681), .A3(new_n624), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NAND4_X1  g504(.A1(new_n681), .A2(new_n640), .A3(new_n475), .A4(new_n592), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  NAND2_X1  g506(.A1(new_n679), .A2(new_n680), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n533), .B1(new_n511), .B2(KEYINPUT70), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n504), .B1(new_n694), .B2(new_n499), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n517), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(G472), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n580), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n571), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n588), .A2(new_n427), .A3(new_n622), .A4(new_n590), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n469), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n693), .A2(new_n701), .A3(new_n575), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  INV_X1    g517(.A(new_n696), .ZN(new_n704));
  INV_X1    g518(.A(new_n698), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n665), .A2(new_n704), .A3(new_n666), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n681), .A2(new_n592), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT105), .B(G125), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G27));
  NAND2_X1  g523(.A1(new_n654), .A2(new_n476), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n317), .B1(new_n678), .B2(new_n295), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n712), .B2(KEYINPUT106), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n714), .B(new_n317), .C1(new_n678), .C2(new_n295), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n714), .B1(new_n313), .B2(new_n317), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n711), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n522), .A2(new_n535), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n584), .B1(new_n722), .B2(new_n518), .ZN(new_n723));
  INV_X1    g537(.A(new_n666), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT42), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n670), .B1(new_n716), .B2(new_n720), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(G131), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G33));
  NAND2_X1  g547(.A1(new_n728), .A2(new_n647), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NAND2_X1  g549(.A1(new_n603), .A2(new_n607), .ZN(new_n736));
  INV_X1    g550(.A(new_n427), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT43), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n583), .A3(new_n632), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n710), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  OAI21_X1  g558(.A(G469), .B1(new_n294), .B2(KEYINPUT45), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n745), .A2(KEYINPUT109), .B1(KEYINPUT45), .B2(new_n294), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n189), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n678), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT110), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n575), .A3(new_n650), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n241), .ZN(G39));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n575), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n754), .B(new_n575), .C1(new_n763), .C2(new_n760), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n538), .A2(new_n571), .A3(new_n666), .A4(new_n710), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT113), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NAND2_X1  g582(.A1(new_n691), .A2(new_n689), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n583), .A2(new_n584), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n623), .A2(KEYINPUT115), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n622), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n427), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n470), .B1(new_n774), .B2(new_n610), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n365), .A2(new_n476), .A3(new_n478), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n770), .A2(new_n777), .A3(new_n712), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n702), .A2(new_n637), .A3(new_n572), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n727), .A2(new_n780), .A3(new_n686), .A4(new_n730), .ZN(new_n781));
  INV_X1    g595(.A(new_n700), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n632), .A2(new_n646), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n659), .A2(new_n782), .A3(new_n712), .A4(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n707), .A2(new_n648), .A3(new_n668), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT52), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n771), .A2(new_n645), .A3(new_n773), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n710), .A2(new_n621), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n640), .A2(new_n789), .A3(new_n712), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n728), .B2(new_n647), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT116), .B1(new_n721), .B2(new_n706), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  INV_X1    g609(.A(new_n706), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n795), .B(new_n796), .C1(new_n716), .C2(new_n720), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n710), .B1(new_n577), .B2(new_n714), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n719), .B1(new_n800), .B2(new_n718), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n715), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n706), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n795), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n721), .A2(KEYINPUT116), .A3(new_n706), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n793), .B1(new_n806), .B2(new_n792), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n787), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n707), .A2(new_n648), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n794), .A2(new_n797), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n734), .A2(new_n790), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n798), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n817), .B2(new_n787), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n808), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n811), .A2(new_n820), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n787), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n693), .B(KEYINPUT114), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n762), .A2(new_n764), .B1(new_n317), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n740), .A2(new_n464), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n699), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n711), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT51), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n655), .A2(new_n476), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n681), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT119), .B1(new_n681), .B2(new_n711), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n644), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n681), .A2(KEYINPUT119), .A3(new_n711), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n659), .A2(new_n584), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n736), .A2(new_n427), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n665), .A2(new_n704), .A3(new_n705), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n839), .A2(new_n844), .A3(new_n740), .A4(new_n840), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n837), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n833), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n832), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n762), .A2(KEYINPUT118), .A3(new_n764), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n828), .A2(new_n317), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n762), .B2(new_n764), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n846), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n847), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n839), .A2(new_n723), .A3(new_n740), .A4(new_n840), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n839), .A2(new_n610), .A3(new_n840), .A4(new_n841), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n681), .A2(new_n592), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n463), .B(G953), .C1(new_n831), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n861), .A2(new_n863), .A3(new_n860), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n826), .A2(new_n870), .B1(G952), .B2(G953), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n873));
  INV_X1    g687(.A(new_n655), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n738), .A2(new_n317), .A3(new_n586), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n841), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n871), .B1(new_n872), .B2(new_n876), .ZN(G75));
  NAND2_X1  g691(.A1(new_n463), .A2(G953), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT122), .Z(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n817), .A2(new_n787), .A3(new_n823), .ZN(new_n881));
  OAI211_X1 g695(.A(G210), .B(G902), .C1(new_n881), .C2(new_n818), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n340), .A2(new_n349), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n348), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT55), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n880), .B1(new_n888), .B2(new_n890), .ZN(G51));
  XNOR2_X1  g705(.A(new_n189), .B(KEYINPUT57), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n881), .A2(new_n818), .A3(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n822), .B1(new_n821), .B2(new_n824), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n675), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n821), .A2(new_n824), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(G902), .A3(new_n746), .A4(new_n747), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n880), .B1(new_n896), .B2(new_n898), .ZN(G54));
  NAND4_X1  g713(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(new_n418), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n418), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n880), .B1(new_n901), .B2(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT59), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n596), .B(new_n905), .C1(new_n893), .C2(new_n894), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n879), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n596), .B1(new_n826), .B2(new_n905), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n897), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n570), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n821), .B2(new_n824), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n880), .B1(new_n916), .B2(new_n630), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n916), .B2(new_n630), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n915), .B(new_n917), .C1(new_n919), .C2(KEYINPUT61), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n630), .B(new_n912), .C1(new_n881), .C2(new_n818), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n879), .C1(new_n916), .C2(new_n570), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n921), .B2(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n467), .B2(new_n346), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT124), .Z(new_n927));
  AND2_X1   g741(.A1(new_n780), .A2(new_n686), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n369), .ZN(new_n930));
  INV_X1    g744(.A(G898), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n885), .B1(new_n931), .B2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n930), .B(new_n932), .ZN(G69));
  XOR2_X1   g747(.A(new_n528), .B(new_n397), .Z(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n642), .B2(new_n369), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n767), .A2(new_n734), .ZN(new_n936));
  INV_X1    g750(.A(new_n731), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n723), .A2(new_n782), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n755), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n809), .A2(new_n668), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n756), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n936), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n935), .B1(new_n942), .B2(new_n369), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n809), .A2(new_n663), .A3(new_n668), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  INV_X1    g759(.A(new_n756), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n711), .B1(new_n774), .B2(new_n610), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n670), .A2(new_n947), .A3(new_n577), .A4(new_n651), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT126), .Z(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n946), .A3(new_n767), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n369), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n934), .B(KEYINPUT125), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n287), .B2(new_n642), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(new_n529), .A2(new_n512), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n936), .A2(new_n941), .A3(new_n937), .A4(new_n928), .ZN(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n950), .A2(new_n929), .ZN(new_n964));
  INV_X1    g778(.A(new_n959), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n656), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n879), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n813), .A2(new_n818), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n529), .A2(new_n499), .ZN(new_n969));
  INV_X1    g783(.A(new_n500), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n959), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n963), .A2(new_n967), .A3(new_n972), .ZN(G57));
endmodule


