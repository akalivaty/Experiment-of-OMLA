//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G125), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AND4_X1   g047(.A1(new_n466), .A2(new_n470), .A3(new_n472), .A4(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n465), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(new_n471), .B2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G137), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n483), .A2(new_n480), .A3(new_n472), .A4(new_n485), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n478), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n475), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G160));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G112), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT72), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  INV_X1    g071(.A(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n483), .A2(new_n480), .A3(new_n497), .A4(new_n472), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n481), .A2(G2105), .A3(new_n483), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n502), .B2(G124), .ZN(G162));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n483), .A2(new_n480), .A3(new_n472), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n497), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT74), .B(G114), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n497), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT4), .A2(G138), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n510), .B(new_n514), .C1(new_n498), .C2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G164));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT75), .B(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  OAI211_X1 g103(.A(G88), .B(new_n519), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(G50), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n531), .B1(new_n529), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND3_X1  g110(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT77), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  OAI21_X1  g118(.A(G543), .B1(new_n527), .B2(new_n528), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT78), .B(G51), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n540), .A2(new_n543), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n520), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n524), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n544), .B1(new_n541), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n523), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n562), .B1(new_n541), .B2(new_n563), .C1(new_n564), .C2(new_n544), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n520), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n542), .A2(G91), .B1(G651), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  OAI21_X1  g157(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n541), .B2(new_n584), .C1(new_n585), .C2(new_n544), .ZN(G288));
  AND2_X1   g161(.A1(new_n519), .A2(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT82), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n524), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(G48), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n541), .C2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n542), .A2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n545), .A2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n523), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G301), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n541), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT83), .ZN(new_n607));
  INV_X1    g182(.A(G651), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n606), .B2(KEYINPUT83), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n545), .A2(G54), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(new_n599), .ZN(G284));
  AOI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(new_n599), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n579), .B(KEYINPUT81), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  XNOR2_X1  g193(.A(G297), .B(KEYINPUT85), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n565), .A2(new_n599), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n620), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g201(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n627));
  NOR3_X1   g202(.A1(new_n471), .A2(new_n469), .A3(G2105), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OAI22_X1  g208(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n631), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n497), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI22_X1  g215(.A1(new_n498), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n502), .B2(G123), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT88), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT90), .Z(new_n664));
  NOR2_X1   g239(.A1(G2072), .A2(G2078), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n443), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(KEYINPUT17), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n667), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n662), .B(new_n663), .C1(new_n443), .C2(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n668), .A3(new_n662), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT91), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NOR2_X1   g269(.A1(G171), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G5), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n694), .A2(G21), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G286), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT99), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT30), .B(G28), .Z(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G29), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n642), .B2(G29), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT98), .Z(new_n709));
  NAND3_X1  g284(.A1(new_n699), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G33), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n497), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n467), .A2(G127), .ZN(new_n715));
  INV_X1    g290(.A(G115), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n469), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n717), .B2(G2105), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n481), .A2(G139), .A3(new_n497), .A4(new_n483), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n712), .B1(new_n720), .B2(new_n711), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G2072), .Z(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n711), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n711), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n728), .A2(new_n729), .B1(G105), .B2(new_n476), .ZN(new_n730));
  INV_X1    g305(.A(G141), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n498), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n502), .B2(G129), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n711), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n711), .B2(G32), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n722), .B1(new_n723), .B2(new_n725), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  OAI22_X1  g315(.A1(G160), .A2(new_n711), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G2084), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n696), .A2(new_n697), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n725), .A2(new_n723), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n745), .B(new_n746), .C1(new_n702), .C2(new_n701), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n710), .A2(new_n737), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n694), .A2(G23), .ZN(new_n750));
  INV_X1    g325(.A(G288), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n694), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT33), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1976), .ZN(new_n754));
  MUX2_X1   g329(.A(G6), .B(G305), .S(G16), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT94), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT32), .B(G1981), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G22), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G166), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1971), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n711), .A2(G25), .ZN(new_n765));
  INV_X1    g340(.A(G131), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n497), .A2(G107), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n498), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n502), .B2(G119), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n765), .B1(new_n775), .B2(new_n711), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT35), .B(G1991), .Z(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n776), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G24), .ZN(new_n780));
  XOR2_X1   g355(.A(G290), .B(KEYINPUT93), .Z(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n763), .A2(new_n764), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n711), .A2(G35), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT102), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n711), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT29), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G2090), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT103), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n694), .A2(G19), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT96), .Z(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n566), .B2(new_n694), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1341), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n711), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT28), .Z(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G116), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n502), .B2(G128), .ZN(new_n804));
  INV_X1    g379(.A(G140), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n498), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n798), .B(new_n811), .C1(G2090), .C2(new_n792), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n694), .A2(G20), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT23), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G299), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  NOR2_X1   g391(.A1(G4), .A2(G16), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n613), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1348), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND4_X1   g395(.A1(new_n794), .A2(new_n812), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n749), .A2(new_n787), .A3(new_n788), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n611), .B(KEYINPUT84), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n620), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n565), .B(KEYINPUT106), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n545), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT105), .B(G93), .Z(new_n832));
  OAI221_X1 g407(.A(new_n830), .B1(new_n523), .B2(new_n831), .C1(new_n541), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n829), .B(new_n833), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT107), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT107), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n824), .B1(KEYINPUT39), .B2(new_n835), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(G145));
  NOR2_X1   g418(.A1(new_n775), .A2(new_n630), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n497), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n498), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n502), .B2(G130), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n774), .A2(new_n629), .ZN(new_n851));
  OR3_X1    g426(.A1(new_n844), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n844), .B2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(new_n720), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n498), .A2(new_n515), .ZN(new_n855));
  INV_X1    g430(.A(G114), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(KEYINPUT74), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(KEYINPUT74), .ZN(new_n858));
  OAI21_X1  g433(.A(G2105), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n859), .A2(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n855), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n808), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n808), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n733), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n865), .A2(new_n733), .A3(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n854), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n720), .A3(new_n867), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n852), .A2(new_n853), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n852), .A2(new_n853), .B1(new_n870), .B2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n873), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G162), .B(new_n490), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n642), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n883), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  INV_X1    g464(.A(KEYINPUT110), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n623), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n623), .A2(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n834), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n829), .B(new_n833), .ZN(new_n895));
  INV_X1    g470(.A(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n617), .A2(KEYINPUT111), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n611), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n617), .A2(KEYINPUT111), .A3(new_n605), .A4(new_n610), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n894), .A2(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n897), .A2(new_n894), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G290), .ZN(new_n912));
  XNOR2_X1  g487(.A(G288), .B(G305), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n912), .B(new_n913), .Z(new_n914));
  INV_X1    g489(.A(new_n910), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n915), .B2(new_n907), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n911), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n833), .A2(new_n599), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(G286), .A2(KEYINPUT112), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(G301), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n924), .B2(G301), .ZN(new_n928));
  NOR2_X1   g503(.A1(G286), .A2(KEYINPUT112), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(G301), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT113), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n933), .B2(new_n926), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n895), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n926), .A3(new_n931), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n834), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n935), .A2(new_n902), .A3(new_n938), .A4(new_n901), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n905), .A2(new_n906), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n935), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(new_n914), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(new_n914), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n923), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n942), .A2(new_n914), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n507), .B2(new_n516), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT67), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n470), .A2(new_n472), .A3(new_n466), .A4(G125), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n464), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G40), .B1(new_n963), .B2(new_n497), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n477), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT115), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n475), .A2(new_n489), .A3(new_n969), .A4(G40), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n958), .B2(KEYINPUT114), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n959), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n808), .B(new_n810), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n733), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT46), .B1(new_n973), .B2(G1996), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n973), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n973), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n733), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT117), .Z(new_n984));
  OAI21_X1  g559(.A(new_n974), .B1(new_n982), .B2(new_n733), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n775), .A2(new_n777), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n774), .A2(new_n778), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT116), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n981), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT48), .Z(new_n994));
  OAI21_X1  g569(.A(new_n980), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n988), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n804), .A2(new_n810), .A3(new_n807), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n973), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n751), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n958), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n964), .A2(new_n967), .A3(KEYINPUT115), .ZN(new_n1003));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n474), .B2(G2105), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n969), .B1(new_n1005), .B2(new_n489), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n958), .B1(new_n968), .B2(new_n970), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT119), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(G305), .A2(G1981), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n1014), .A2(new_n1015), .A3(KEYINPUT49), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT49), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT121), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1015), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1009), .A2(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n1001), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1013), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(new_n1000), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT120), .B(G1976), .Z(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1027), .A2(new_n1029), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n1031), .B2(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT55), .Z(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n958), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT45), .B(new_n957), .C1(new_n507), .C2(new_n516), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n971), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT118), .B(G1971), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n863), .A2(new_n1042), .A3(new_n957), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2090), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n971), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1011), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1025), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1025), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1034), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1055), .A2(new_n1056), .A3(G2090), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1039), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1037), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n863), .B2(new_n957), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1061), .B2(new_n971), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1030), .A2(new_n1032), .A3(new_n1054), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G286), .A2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n702), .B1(new_n1055), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2084), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n971), .A2(new_n1070), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1966), .B1(new_n1061), .B2(new_n971), .ZN(new_n1074));
  OAI21_X1  g649(.A(G8), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1067), .B2(KEYINPUT123), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1067), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1080));
  OAI211_X1 g655(.A(G8), .B(new_n1077), .C1(new_n1080), .C2(G286), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1038), .B2(G2078), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n697), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1061), .A2(KEYINPUT53), .A3(new_n723), .A4(new_n971), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n497), .B1(new_n474), .B2(KEYINPUT124), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(KEYINPUT124), .B2(new_n474), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1083), .A2(new_n1004), .A3(G2078), .ZN(new_n1093));
  AND4_X1   g668(.A1(new_n489), .A2(new_n1092), .A3(new_n1037), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n959), .A2(new_n972), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1088), .A2(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n1085), .A3(new_n1084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1066), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1007), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1061), .A2(new_n982), .A3(new_n971), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n1103), .B2(new_n566), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1105), .B(new_n565), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n819), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1010), .A2(new_n810), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n825), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n613), .A2(new_n1108), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n574), .A2(new_n1117), .A3(new_n578), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n574), .B2(new_n578), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1061), .A2(new_n971), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1120), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1122), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1107), .A2(new_n1116), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n825), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1125), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1054), .A2(new_n1065), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1075), .A2(G286), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1032), .A3(new_n1030), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1099), .A2(new_n1135), .B1(KEYINPUT63), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1082), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1087), .A2(G171), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1066), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n1082), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1082), .A2(new_n1145), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1138), .A2(KEYINPUT63), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1053), .A2(new_n1139), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  AND2_X1   g726(.A1(G290), .A2(G1986), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n992), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n990), .B1(new_n981), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n999), .B1(new_n1155), .B2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g732(.A1(G401), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1159));
  INV_X1    g733(.A(new_n886), .ZN(new_n1160));
  AOI21_X1  g734(.A(new_n884), .B1(new_n878), .B2(new_n879), .ZN(new_n1161));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n1162), .B1(new_n953), .B2(new_n954), .ZN(G308));
  OAI221_X1 g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1160), .C1(new_n947), .C2(new_n948), .ZN(G225));
endmodule


