//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT66), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G107), .C2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n212), .B(new_n232), .C1(new_n235), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G238), .B(G244), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(G107), .ZN(new_n249));
  INV_X1    g0049(.A(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n202), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT69), .B(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(G274), .C1(new_n259), .C2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n229), .A2(G1698), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(G226), .C2(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n260), .B1(new_n214), .B2(new_n265), .C1(new_n270), .C2(new_n263), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n271), .A2(new_n272), .ZN(new_n274));
  OAI21_X1  g0074(.A(G169), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT14), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT77), .ZN(new_n278));
  INV_X1    g0078(.A(new_n274), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT77), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n271), .A2(new_n280), .A3(KEYINPUT13), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(G179), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n271), .B(new_n272), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G169), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n276), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n234), .A3(G1), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT79), .B1(new_n289), .B2(G68), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT12), .Z(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n233), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G1), .B2(new_n234), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n291), .B1(new_n213), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n261), .A2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G77), .B1(G20), .B2(new_n213), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n234), .A2(new_n261), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n202), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n293), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n286), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n283), .A2(G200), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n307), .B(new_n304), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT80), .Z(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n288), .A2(G50), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n295), .B2(G50), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n204), .A2(G20), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n299), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n319), .A2(new_n297), .B1(G150), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n294), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n323), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT74), .B1(new_n323), .B2(KEYINPUT9), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G222), .ZN(new_n328));
  INV_X1    g0128(.A(G223), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n266), .B(new_n328), .C1(new_n329), .C2(new_n327), .ZN(new_n330));
  INV_X1    g0130(.A(new_n263), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(G77), .C2(new_n266), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n260), .C1(new_n224), .C2(new_n265), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(new_n309), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(KEYINPUT9), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n326), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT10), .ZN(new_n338));
  INV_X1    g0138(.A(new_n323), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n333), .A2(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n329), .A2(new_n327), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n224), .A2(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n266), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n331), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n265), .A2(new_n229), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n260), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT83), .B1(new_n353), .B2(G190), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n263), .B1(new_n347), .B2(new_n348), .ZN(new_n357));
  INV_X1    g0157(.A(new_n260), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(new_n358), .A3(new_n351), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT83), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n309), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n366), .B2(new_n234), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n368), .B(G20), .C1(new_n363), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n299), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n234), .B1(new_n236), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n368), .B1(new_n266), .B2(G20), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n364), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT7), .B(new_n234), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n375), .B1(new_n384), .B2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n373), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n293), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n318), .A2(new_n288), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n295), .B2(new_n318), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n362), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT82), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n353), .A2(new_n340), .ZN(new_n395));
  INV_X1    g0195(.A(G179), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n350), .A2(new_n396), .A3(new_n352), .A4(new_n260), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n385), .B2(new_n373), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n213), .B1(new_n380), .B2(new_n383), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n400), .A2(new_n378), .A3(new_n372), .A4(new_n375), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n399), .A2(new_n401), .A3(new_n294), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(new_n389), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n394), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n395), .A2(new_n397), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n387), .B2(new_n390), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n407), .A2(KEYINPUT82), .A3(KEYINPUT18), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n387), .A2(new_n390), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT18), .A4(new_n398), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n407), .B2(KEYINPUT18), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n393), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n287), .A2(G20), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n258), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n258), .B2(new_n234), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n225), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n297), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT71), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n299), .B2(new_n318), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(new_n423), .B2(new_n293), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n288), .A2(new_n225), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n425), .B(KEYINPUT72), .Z(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G238), .A2(G1698), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n266), .B(new_n428), .C1(new_n229), .C2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n331), .C1(G107), .C2(new_n266), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n260), .C1(new_n226), .C2(new_n265), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n340), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT73), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n431), .A2(G179), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(KEYINPUT73), .A3(new_n432), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n431), .A2(new_n309), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(G200), .B2(new_n431), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(new_n424), .A3(new_n426), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n415), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n312), .A2(new_n344), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n289), .B(new_n294), .C1(G1), .C2(new_n261), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT25), .B1(new_n288), .B2(new_n445), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n444), .A2(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT90), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n363), .A2(new_n365), .A3(new_n234), .A4(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n266), .A2(new_n454), .A3(new_n234), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n261), .A2(new_n250), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n234), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n234), .A2(G107), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT23), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n453), .A2(new_n455), .B1(new_n234), .B2(new_n457), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n451), .B1(new_n466), .B2(new_n293), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT90), .B(new_n294), .C1(new_n462), .C2(new_n465), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n450), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n363), .A2(new_n365), .A3(G257), .A4(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT91), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n266), .A2(new_n472), .A3(G257), .A4(G1698), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT93), .B(G294), .Z(new_n474));
  OAI211_X1 g0274(.A(new_n471), .B(new_n473), .C1(new_n261), .C2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n266), .A2(G250), .A3(new_n327), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT92), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n266), .A2(KEYINPUT92), .A3(G250), .A4(new_n327), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n331), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n263), .A2(G274), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n259), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n258), .A2(G45), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT86), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n490), .B(new_n487), .C1(new_n259), .C2(new_n485), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n484), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n487), .B1(new_n259), .B2(new_n485), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n331), .B1(new_n493), .B2(new_n482), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G264), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n481), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT94), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(KEYINPUT94), .A3(G264), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n481), .A2(new_n499), .A3(new_n492), .A4(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n497), .A2(new_n309), .B1(new_n501), .B2(new_n355), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n469), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n464), .B1(new_n463), .B2(new_n460), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n293), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n466), .A2(new_n451), .A3(new_n293), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n449), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n492), .A2(new_n481), .A3(new_n499), .A4(new_n500), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(G179), .B1(G169), .B2(new_n496), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT95), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT95), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n497), .A2(new_n340), .B1(new_n501), .B2(new_n396), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n469), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n503), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n288), .A2(new_n250), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n234), .C1(G33), .C2(new_n218), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n293), .C1(new_n234), .C2(G116), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT20), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n517), .B1(new_n250), .B2(new_n444), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n494), .A2(G270), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G264), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n266), .B(new_n527), .C1(new_n219), .C2(G1698), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n331), .C1(G303), .C2(new_n266), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n492), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n525), .A2(new_n396), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n524), .A2(new_n530), .A3(G169), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(G200), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n525), .C1(new_n309), .C2(new_n530), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n363), .A2(new_n365), .A3(G244), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n540), .A2(new_n541), .B1(G33), .B2(G283), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n327), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n266), .A2(G250), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n327), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT85), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n366), .A2(new_n217), .ZN(new_n548));
  OAI21_X1  g0348(.A(G1698), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n542), .A4(new_n543), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n551), .A3(new_n331), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n494), .A2(G257), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n492), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n554), .A3(G190), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n299), .A2(new_n225), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n218), .A2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g0359(.A(G97), .B(G107), .Z(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n561), .B2(G20), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n384), .A2(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n294), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n444), .A2(new_n218), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n289), .A2(G97), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n555), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n355), .B1(new_n552), .B2(new_n554), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n539), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n552), .A2(new_n554), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(KEYINPUT87), .A3(new_n567), .A4(new_n555), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n567), .B1(new_n340), .B2(new_n571), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n552), .A2(new_n554), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(KEYINPUT88), .A3(new_n396), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT88), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n571), .B2(G179), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n487), .A2(new_n217), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n263), .B(new_n581), .C1(G274), .C2(new_n487), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G238), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n226), .B2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n457), .B1(new_n584), .B2(new_n266), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n582), .B1(new_n585), .B2(new_n263), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G169), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n396), .B2(new_n586), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT89), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n266), .A2(new_n234), .A3(G68), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n216), .A2(new_n218), .A3(new_n445), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n269), .A2(new_n234), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT19), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n269), .A2(G20), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n590), .B(new_n593), .C1(KEYINPUT19), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n420), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n293), .B1(new_n288), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n596), .B2(new_n444), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n586), .A2(new_n309), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n586), .A2(G200), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n444), .A2(new_n216), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n589), .A2(new_n598), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n574), .A2(new_n580), .A3(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n443), .A2(new_n516), .A3(new_n538), .A4(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n588), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n602), .A2(new_n599), .B1(new_n598), .B2(new_n588), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n575), .A2(new_n577), .A3(new_n579), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n603), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT26), .B1(new_n612), .B2(new_n580), .ZN(new_n613));
  INV_X1    g0413(.A(new_n608), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n510), .A2(G200), .B1(G190), .B2(new_n496), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n509), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n535), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n509), .A2(new_n511), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n574), .A2(new_n580), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n611), .B(new_n613), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n443), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n343), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n310), .B1(new_n305), .B2(new_n286), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT18), .B(new_n398), .C1(new_n402), .C2(new_n389), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n407), .A2(KEYINPUT18), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n625), .A2(new_n393), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n629), .B2(new_n338), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n622), .A2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n258), .A2(new_n234), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n618), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  INV_X1    g0439(.A(new_n637), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n516), .B1(new_n509), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n535), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n618), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n642), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n524), .A2(new_n637), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n538), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n535), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n647), .A2(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n259), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n209), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n591), .A2(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n237), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n604), .A2(new_n516), .A3(new_n538), .A4(new_n640), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n586), .A2(new_n396), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n481), .A2(new_n499), .A3(new_n500), .A4(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n492), .A2(new_n526), .A3(new_n529), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n576), .A2(new_n664), .A3(KEYINPUT30), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(G179), .B1(new_n552), .B2(new_n554), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n501), .A3(new_n530), .A4(new_n586), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n552), .A3(new_n554), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n481), .A2(new_n499), .A3(new_n500), .A4(new_n663), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n666), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT31), .B1(new_n673), .B2(new_n637), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT97), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n637), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT97), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n674), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n662), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT98), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(KEYINPUT98), .A3(G330), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n621), .A2(new_n640), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n512), .A2(new_n515), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n535), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT99), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n574), .A2(new_n694), .A3(new_n580), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n574), .B2(new_n580), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n693), .B(new_n616), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n612), .A2(new_n580), .A3(KEYINPUT26), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .A3(new_n640), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n689), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n661), .B1(new_n705), .B2(G1), .ZN(G364));
  NAND3_X1  g0506(.A1(G355), .A2(new_n209), .A3(new_n266), .ZN(new_n707));
  INV_X1    g0507(.A(G45), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n256), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n366), .A2(new_n209), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G45), .B2(new_n237), .ZN(new_n712));
  OAI221_X1 g0512(.A(new_n707), .B1(G116), .B2(new_n209), .C1(new_n709), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n233), .B1(G20), .B2(new_n340), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT101), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n234), .A2(new_n309), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n355), .A2(G179), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n216), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n396), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n396), .A2(new_n355), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n266), .B1(new_n726), .B2(new_n228), .C1(new_n202), .C2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n234), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n371), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT32), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n722), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n734), .B1(new_n445), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G97), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n727), .A2(new_n730), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n213), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n729), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n725), .A2(new_n730), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n225), .B2(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n724), .B(new_n744), .C1(new_n734), .C2(new_n733), .ZN(new_n745));
  INV_X1    g0545(.A(new_n740), .ZN(new_n746));
  INV_X1    g0546(.A(G317), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT33), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(KEYINPUT33), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n732), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n750), .B(new_n752), .C1(new_n753), .C2(new_n735), .ZN(new_n754));
  INV_X1    g0554(.A(new_n728), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(G326), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n474), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n738), .ZN(new_n758));
  INV_X1    g0558(.A(new_n723), .ZN(new_n759));
  INV_X1    g0559(.A(new_n726), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G303), .A2(new_n759), .B1(new_n760), .B2(G322), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n756), .A2(new_n366), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n743), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G311), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n745), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT102), .Z(new_n766));
  AOI21_X1  g0566(.A(new_n720), .B1(new_n766), .B2(new_n717), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n416), .A2(G45), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n657), .A2(G1), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n716), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n767), .B(new_n770), .C1(new_n651), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n651), .A2(G330), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n652), .A2(new_n769), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(G396));
  NAND2_X1  g0575(.A1(new_n427), .A2(new_n637), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n438), .A2(new_n441), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n438), .B2(new_n776), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n621), .A2(new_n640), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n778), .B(KEYINPUT104), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n690), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n688), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n769), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n739), .B1(new_n445), .B2(new_n723), .C1(new_n784), .C2(new_n732), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n366), .B1(new_n726), .B2(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n216), .A2(new_n735), .B1(new_n743), .B2(new_n250), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n753), .B2(new_n740), .C1(new_n790), .C2(new_n728), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n732), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G143), .A2(new_n760), .B1(new_n763), .B2(G159), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n755), .A2(G137), .ZN(new_n795));
  INV_X1    g0595(.A(G150), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n740), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  AOI211_X1 g0598(.A(new_n793), .B(new_n798), .C1(G50), .C2(new_n759), .ZN(new_n799));
  INV_X1    g0599(.A(new_n738), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n228), .B2(new_n800), .C1(new_n213), .C2(new_n735), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n791), .B1(new_n801), .B2(new_n366), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n769), .B1(new_n802), .B2(new_n717), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n717), .A2(new_n714), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(G77), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT103), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n715), .B2(new_n778), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n783), .A2(new_n808), .ZN(G384));
  AOI21_X1  g0609(.A(new_n250), .B1(new_n561), .B2(KEYINPUT35), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n810), .B(new_n235), .C1(KEYINPUT35), .C2(new_n561), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT36), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n374), .A2(G77), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n237), .A2(new_n813), .B1(G50), .B2(new_n213), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(G1), .A3(new_n287), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n305), .A2(new_n637), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n306), .A2(new_n310), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n286), .A2(new_n305), .A3(new_n637), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n778), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT108), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n674), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n680), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n678), .A2(new_n821), .A3(new_n679), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n662), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT105), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n635), .B1(new_n387), .B2(new_n390), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n828), .B1(new_n415), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n403), .A3(new_n391), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n403), .A2(new_n394), .A3(new_n404), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n626), .A2(KEYINPUT81), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT82), .B1(new_n407), .B2(KEYINPUT18), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT18), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n391), .B(KEYINPUT17), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(KEYINPUT105), .A3(new_n829), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n831), .A2(KEYINPUT38), .A3(new_n833), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n627), .A2(new_n628), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n829), .B1(new_n393), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n832), .A2(KEYINPUT106), .A3(KEYINPUT37), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(new_n833), .C2(KEYINPUT106), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n827), .A2(new_n849), .A3(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(new_n662), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n778), .B(new_n819), .C1(new_n851), .C2(new_n825), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n831), .A2(new_n833), .A3(new_n841), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n847), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n852), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n855), .A2(KEYINPUT109), .A3(KEYINPUT40), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT109), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT105), .B1(new_n840), .B2(new_n829), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n828), .B(new_n830), .C1(new_n838), .C2(new_n839), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n860), .B2(new_n833), .ZN(new_n861));
  AND4_X1   g0661(.A1(KEYINPUT38), .A2(new_n831), .A3(new_n833), .A4(new_n841), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n827), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(G330), .B(new_n850), .C1(new_n856), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n851), .A2(new_n825), .ZN(new_n867));
  INV_X1    g0667(.A(G330), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n443), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n850), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT109), .B1(new_n855), .B2(KEYINPUT40), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n863), .A2(new_n857), .A3(new_n864), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n851), .B2(new_n825), .ZN(new_n876));
  INV_X1    g0676(.A(new_n443), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n842), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n849), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n306), .A2(new_n637), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n854), .A2(new_n842), .ZN(new_n884));
  INV_X1    g0684(.A(new_n819), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n624), .A2(new_n640), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n779), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n884), .A2(new_n887), .B1(new_n843), .B2(new_n635), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT107), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n883), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n878), .B(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n443), .A2(new_n691), .A3(new_n702), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n630), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n812), .B(new_n815), .C1(new_n896), .C2(new_n417), .ZN(G367));
  NOR2_X1   g0697(.A1(new_n695), .A2(new_n696), .ZN(new_n898));
  INV_X1    g0698(.A(new_n567), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n637), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n580), .A2(new_n640), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n654), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n644), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n640), .B1(new_n597), .B2(new_n601), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n607), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n614), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n512), .A3(new_n515), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n580), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(KEYINPUT110), .A3(new_n580), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n640), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n905), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT111), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n909), .B1(new_n905), .B2(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n903), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n768), .A2(G1), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n643), .B1(new_n651), .B2(G330), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n648), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n704), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n646), .A2(new_n902), .A3(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n646), .A2(new_n902), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT112), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT44), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT45), .B1(new_n646), .B2(new_n902), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n646), .A2(new_n902), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n705), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n657), .B(KEYINPUT41), .Z(new_n938));
  AOI21_X1  g0738(.A(new_n924), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n918), .A2(new_n903), .A3(new_n921), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n923), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n800), .A2(new_n213), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n266), .B1(new_n735), .B2(new_n225), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT113), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n760), .A2(G150), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G143), .A2(new_n755), .B1(new_n759), .B2(G58), .ZN(new_n947));
  AOI22_X1  g0747(.A1(G50), .A2(new_n763), .B1(new_n751), .B2(G137), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n943), .B(new_n949), .C1(G159), .C2(new_n746), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n738), .A2(G107), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G303), .A2(new_n760), .B1(new_n751), .B2(G317), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n366), .C1(new_n218), .C2(new_n735), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n757), .A2(new_n746), .B1(new_n763), .B2(G283), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n784), .B2(new_n728), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n723), .A2(new_n250), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n950), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n717), .ZN(new_n961));
  INV_X1    g0761(.A(new_n711), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n719), .B1(new_n209), .B2(new_n596), .C1(new_n242), .C2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n908), .A2(new_n771), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n961), .A2(new_n770), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n942), .A2(new_n965), .ZN(G387));
  NAND2_X1  g0766(.A1(new_n648), .A2(new_n716), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n318), .A2(KEYINPUT50), .A3(G50), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT50), .B1(new_n318), .B2(G50), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n708), .A4(new_n658), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n213), .A2(new_n225), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n711), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT114), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n708), .B2(new_n247), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n266), .A2(new_n209), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(G107), .B2(new_n209), .C1(new_n658), .C2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n719), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n759), .A2(G77), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n371), .B2(new_n728), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n800), .A2(new_n596), .B1(new_n726), .B2(new_n202), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n751), .A2(G150), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n366), .B1(new_n746), .B2(new_n319), .ZN(new_n984));
  INV_X1    g0784(.A(new_n735), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G68), .A2(new_n763), .B1(new_n985), .B2(G97), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G322), .A2(new_n755), .B1(new_n746), .B2(G311), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n790), .B2(new_n743), .C1(new_n747), .C2(new_n726), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n753), .B2(new_n800), .C1(new_n474), .C2(new_n723), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT49), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n266), .B1(new_n751), .B2(G326), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n250), .B2(new_n735), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n987), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n717), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n967), .A2(new_n770), .A3(new_n978), .A4(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n924), .ZN(new_n998));
  INV_X1    g0798(.A(new_n657), .ZN(new_n999));
  INV_X1    g0799(.A(new_n926), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n705), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n997), .B1(new_n998), .B2(new_n926), .C1(new_n1001), .C2(new_n927), .ZN(G393));
  INV_X1    g0802(.A(KEYINPUT116), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n935), .B1(new_n1003), .B2(new_n653), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n654), .A2(KEYINPUT116), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n999), .B(new_n936), .C1(new_n1006), .C2(new_n927), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n728), .A2(new_n747), .B1(new_n726), .B2(new_n784), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT52), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G116), .B2(new_n738), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n445), .A2(new_n735), .B1(new_n743), .B2(new_n786), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n266), .B(new_n1011), .C1(G322), .C2(new_n751), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n790), .C2(new_n740), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G283), .B2(new_n759), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n740), .A2(new_n202), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n723), .A2(new_n213), .B1(new_n743), .B2(new_n318), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G77), .C2(new_n738), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G87), .A2(new_n985), .B1(new_n751), .B2(G143), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n728), .A2(new_n796), .B1(new_n726), .B2(new_n371), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  AND4_X1   g0820(.A1(new_n266), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n717), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n719), .B1(new_n218), .B2(new_n209), .C1(new_n253), .C2(new_n962), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT117), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n770), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n902), .B2(new_n716), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1006), .B2(new_n924), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1007), .A2(new_n1027), .ZN(G390));
  NOR3_X1   g0828(.A1(new_n867), .A2(new_n868), .A3(new_n820), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n779), .A2(new_n886), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n882), .B1(new_n1030), .B2(new_n819), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n879), .B2(new_n881), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n701), .A2(new_n640), .A3(new_n778), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n885), .B1(new_n1033), .B2(new_n886), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n882), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n849), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1029), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n688), .A2(new_n778), .A3(new_n819), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT118), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n1029), .C1(new_n1032), .C2(new_n1037), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1039), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1033), .A2(new_n886), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n869), .A2(new_n780), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n885), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1041), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n687), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT98), .B1(new_n683), .B2(G330), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n778), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1029), .B1(new_n1052), .B2(new_n885), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1030), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n894), .A2(new_n630), .A3(new_n870), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1045), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n819), .B1(new_n688), .B2(new_n778), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1030), .B1(new_n1060), .B2(new_n1029), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1056), .B1(new_n1061), .B2(new_n1049), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1062), .A2(new_n1042), .A3(new_n1044), .A4(new_n1039), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1063), .A3(new_n999), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1045), .A2(new_n998), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n879), .A2(new_n881), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n714), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n804), .A2(new_n318), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(new_n743), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n759), .A2(G150), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT53), .ZN(new_n1073));
  INV_X1    g0873(.A(G125), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n266), .B1(new_n732), .B2(new_n1074), .C1(new_n792), .C2(new_n726), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n755), .A2(G128), .B1(new_n985), .B2(G50), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n371), .C2(new_n800), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1071), .B(new_n1078), .C1(G137), .C2(new_n746), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n728), .A2(new_n753), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n724), .B1(G68), .B2(new_n985), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n746), .A2(G107), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n266), .B1(new_n738), .B2(G77), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G97), .A2(new_n763), .B1(new_n751), .B2(G294), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1080), .B(new_n1085), .C1(G116), .C2(new_n760), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n717), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1067), .A2(new_n770), .A3(new_n1068), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1064), .A2(new_n1065), .A3(new_n1088), .ZN(G378));
  OAI221_X1 g0889(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n259), .C2(new_n266), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n979), .B1(new_n732), .B2(new_n753), .C1(new_n250), .C2(new_n728), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n746), .A2(G97), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n760), .A2(G107), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n985), .A2(G58), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n259), .A2(new_n266), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n596), .A2(new_n743), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1091), .A2(new_n1096), .A3(new_n943), .A4(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT58), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n1069), .A2(new_n759), .B1(new_n760), .B2(G128), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT119), .Z(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n1074), .B2(new_n728), .C1(new_n792), .C2(new_n740), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G137), .B2(new_n763), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n796), .B2(new_n800), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT59), .ZN(new_n1105));
  AOI211_X1 g0905(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n371), .B2(new_n735), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1090), .B(new_n1099), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n769), .B1(new_n1108), .B2(new_n717), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n344), .B(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n323), .A2(new_n635), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n344), .B(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1109), .B1(G50), .B2(new_n805), .C1(new_n1119), .C2(new_n715), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n890), .A2(new_n891), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n873), .A2(new_n874), .ZN(new_n1122));
  AND4_X1   g0922(.A1(G330), .A2(new_n1122), .A3(new_n850), .A4(new_n1118), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1118), .B1(new_n875), .B2(G330), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n866), .A2(new_n1119), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n875), .A2(G330), .A3(new_n1118), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n892), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n998), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1125), .A2(new_n1128), .B1(new_n1063), .B2(new_n1057), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n999), .B1(new_n1131), .B2(KEYINPUT57), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT120), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1125), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1063), .B2(new_n1057), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1126), .A2(new_n892), .A3(new_n1127), .A4(KEYINPUT120), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1120), .B(new_n1130), .C1(new_n1132), .C2(new_n1138), .ZN(G375));
  NAND3_X1  g0939(.A1(new_n1061), .A2(new_n1056), .A3(new_n1049), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n938), .B(KEYINPUT121), .Z(new_n1141));
  NAND3_X1  g0941(.A1(new_n1058), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n723), .A2(new_n218), .B1(new_n735), .B2(new_n225), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n800), .A2(new_n596), .B1(new_n790), .B2(new_n732), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G294), .C2(new_n755), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n266), .B1(new_n763), .B2(G107), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n753), .C2(new_n726), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G116), .B2(new_n746), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1094), .B1(new_n792), .B2(new_n728), .C1(new_n202), .C2(new_n800), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G137), .B2(new_n760), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n751), .A2(G128), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n266), .B1(new_n743), .B2(new_n796), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G159), .B2(new_n759), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n746), .B2(new_n1069), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n717), .B1(new_n1148), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n770), .B(new_n1156), .C1(new_n819), .C2(new_n715), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n213), .B2(new_n804), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1055), .B2(new_n924), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1142), .A2(new_n1159), .ZN(G381));
  OAI21_X1  g0960(.A(new_n1057), .B1(new_n1045), .B2(new_n1058), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1126), .A2(new_n892), .A3(new_n1127), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n892), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n657), .B1(new_n1164), .B2(new_n1135), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1129), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(G378), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n1120), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n942), .A2(new_n965), .A3(new_n1027), .A4(new_n1007), .ZN(new_n1170));
  OR3_X1    g0970(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1170), .A2(G384), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1169), .B1(new_n1172), .B2(KEYINPUT122), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT122), .B2(new_n1172), .ZN(G407));
  OAI211_X1 g0974(.A(G407), .B(G213), .C1(G343), .C2(new_n1169), .ZN(G409));
  NAND2_X1  g0975(.A1(G375), .A2(G378), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1134), .A2(new_n924), .A3(new_n1137), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1120), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT123), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT123), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1180), .A3(new_n1120), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1168), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n636), .A2(G213), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT125), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1140), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1061), .A2(KEYINPUT60), .A3(new_n1056), .A4(new_n1049), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n999), .A3(new_n1058), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1159), .ZN(new_n1190));
  INV_X1    g0990(.A(G384), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1185), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(KEYINPUT125), .B(G384), .C1(new_n1189), .C2(new_n1159), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1189), .A2(G384), .A3(new_n1159), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT124), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT124), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1189), .A2(new_n1198), .A3(G384), .A4(new_n1159), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1193), .A2(new_n1195), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1176), .A2(new_n1183), .A3(new_n1184), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT62), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1176), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1184), .A2(KEYINPUT126), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1207), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1204), .A3(new_n1210), .A4(new_n1205), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1203), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G375), .A2(G378), .B1(G213), .B2(new_n636), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT62), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1183), .A4(new_n1200), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1202), .A2(new_n1213), .A3(new_n1214), .A4(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n918), .A2(new_n903), .A3(new_n921), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(new_n922), .A3(new_n939), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n965), .ZN(new_n1221));
  OAI21_X1  g1021(.A(G390), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(G393), .B(G396), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1222), .A2(new_n1170), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1222), .B2(new_n1170), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1218), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1215), .A2(KEYINPUT63), .A3(new_n1183), .A4(new_n1200), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1229), .A2(new_n1214), .A3(new_n1226), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1215), .A2(new_n1183), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT63), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1201), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(G405));
  NAND2_X1  g1035(.A1(new_n1209), .A2(new_n1204), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1176), .A2(new_n1169), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1176), .B2(new_n1169), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1237), .A2(new_n1238), .A3(KEYINPUT127), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G375), .A2(G378), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1168), .B1(new_n1167), .B2(new_n1120), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1200), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1176), .A2(new_n1169), .A3(new_n1236), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1227), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT127), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1226), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(G402));
endmodule


