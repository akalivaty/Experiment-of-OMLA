

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  NOR2_X1 U323 ( .A1(n473), .A2(n575), .ZN(n475) );
  INV_X1 U324 ( .A(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U325 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n431) );
  XNOR2_X1 U327 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U328 ( .A(n454), .B(KEYINPUT121), .ZN(n571) );
  XOR2_X1 U329 ( .A(KEYINPUT28), .B(n466), .Z(n542) );
  XNOR2_X1 U330 ( .A(n343), .B(n342), .ZN(n528) );
  XNOR2_X1 U331 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U332 ( .A(G92GAT), .B(G85GAT), .Z(n291) );
  NAND2_X1 U333 ( .A1(n328), .A2(n466), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U335 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n459) );
  INV_X1 U336 ( .A(KEYINPUT93), .ZN(n334) );
  XNOR2_X1 U337 ( .A(n528), .B(n459), .ZN(n468) );
  INV_X1 U338 ( .A(KEYINPUT104), .ZN(n478) );
  INV_X1 U339 ( .A(KEYINPUT19), .ZN(n330) );
  XNOR2_X1 U340 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U341 ( .A(n433), .B(KEYINPUT54), .ZN(n434) );
  XNOR2_X1 U342 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U343 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U344 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U345 ( .A(n333), .B(n332), .ZN(n450) );
  XNOR2_X1 U346 ( .A(n402), .B(n401), .ZN(n426) );
  XNOR2_X1 U347 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U348 ( .A(n426), .B(KEYINPUT41), .ZN(n558) );
  INV_X1 U349 ( .A(G29GAT), .ZN(n485) );
  XNOR2_X1 U350 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n483) );
  XNOR2_X1 U352 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U353 ( .A(n484), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U354 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n294) );
  XNOR2_X1 U355 ( .A(KEYINPUT1), .B(KEYINPUT90), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U357 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n295) );
  XOR2_X1 U358 ( .A(n295), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U359 ( .A(G162GAT), .B(n314), .ZN(n297) );
  XOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .Z(n449) );
  XNOR2_X1 U361 ( .A(G134GAT), .B(n449), .ZN(n296) );
  XNOR2_X1 U362 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n312) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G120GAT), .Z(n301) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U366 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U367 ( .A(G57GAT), .B(G148GAT), .Z(n303) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G141GAT), .ZN(n302) );
  XNOR2_X1 U369 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U370 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U371 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n307) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U374 ( .A(KEYINPUT92), .B(n308), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n575) );
  INV_X1 U377 ( .A(n575), .ZN(n328) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n313), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U380 ( .A(n337), .B(n314), .ZN(n327) );
  XOR2_X1 U381 ( .A(G50GAT), .B(G162GAT), .Z(n417) );
  XOR2_X1 U382 ( .A(G148GAT), .B(G78GAT), .Z(n386) );
  XOR2_X1 U383 ( .A(n417), .B(n386), .Z(n316) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U385 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U386 ( .A(KEYINPUT22), .B(G204GAT), .Z(n318) );
  XNOR2_X1 U387 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n317) );
  XNOR2_X1 U388 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U389 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U390 ( .A(G141GAT), .B(G22GAT), .Z(n367) );
  XOR2_X1 U391 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n322) );
  XNOR2_X1 U392 ( .A(G218GAT), .B(G106GAT), .ZN(n321) );
  XNOR2_X1 U393 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U394 ( .A(n367), .B(n323), .ZN(n324) );
  XNOR2_X1 U395 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n466) );
  XNOR2_X1 U397 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n329) );
  XNOR2_X1 U398 ( .A(n329), .B(KEYINPUT18), .ZN(n333) );
  XNOR2_X1 U399 ( .A(G169GAT), .B(G176GAT), .ZN(n331) );
  XNOR2_X1 U400 ( .A(n450), .B(G190GAT), .ZN(n341) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U402 ( .A(G204GAT), .B(G64GAT), .Z(n398) );
  XOR2_X1 U403 ( .A(n398), .B(G92GAT), .Z(n338) );
  XOR2_X1 U404 ( .A(G36GAT), .B(G218GAT), .Z(n415) );
  XOR2_X1 U405 ( .A(G8GAT), .B(KEYINPUT78), .Z(n357) );
  XOR2_X1 U406 ( .A(n415), .B(n357), .Z(n342) );
  XOR2_X1 U407 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n345) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n363) );
  XOR2_X1 U410 ( .A(G211GAT), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U413 ( .A(G64GAT), .B(G78GAT), .Z(n349) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(G155GAT), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U416 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U417 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n353) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U420 ( .A(KEYINPUT82), .B(n354), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U422 ( .A(n358), .B(n357), .Z(n361) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G127GAT), .Z(n444) );
  XNOR2_X1 U424 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n359), .B(KEYINPUT71), .ZN(n387) );
  XNOR2_X1 U426 ( .A(n444), .B(n387), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n570) );
  XOR2_X1 U429 ( .A(G15GAT), .B(G113GAT), .Z(n365) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(G50GAT), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U432 ( .A(n366), .B(G36GAT), .Z(n369) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(n367), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U435 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT7), .ZN(n418) );
  XOR2_X1 U437 ( .A(n418), .B(KEYINPUT68), .Z(n372) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U440 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT30), .B(G8GAT), .Z(n376) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G1GAT), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U444 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n378) );
  XNOR2_X1 U445 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n568) );
  XNOR2_X1 U449 ( .A(G99GAT), .B(G106GAT), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n291), .B(n383), .ZN(n412) );
  XNOR2_X1 U451 ( .A(n412), .B(KEYINPUT33), .ZN(n385) );
  AND2_X1 U452 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U454 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XOR2_X1 U455 ( .A(n443), .B(n386), .Z(n388) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n393) );
  INV_X1 U457 ( .A(n393), .ZN(n391) );
  NAND2_X1 U458 ( .A1(n391), .A2(KEYINPUT72), .ZN(n395) );
  INV_X1 U459 ( .A(KEYINPUT72), .ZN(n392) );
  NAND2_X1 U460 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U461 ( .A1(n395), .A2(n394), .ZN(n402) );
  XOR2_X1 U462 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n397) );
  XNOR2_X1 U463 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n396) );
  XOR2_X1 U464 ( .A(n397), .B(n396), .Z(n400) );
  XNOR2_X1 U465 ( .A(G176GAT), .B(n398), .ZN(n399) );
  AND2_X1 U466 ( .A1(n568), .A2(n558), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(KEYINPUT46), .ZN(n404) );
  NOR2_X1 U468 ( .A1(n570), .A2(n404), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT112), .ZN(n423) );
  XOR2_X1 U470 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT66), .B(KEYINPUT11), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n422) );
  XOR2_X1 U473 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n409) );
  NAND2_X1 U474 ( .A1(G232GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U476 ( .A(n410), .B(KEYINPUT75), .Z(n414) );
  XNOR2_X1 U477 ( .A(G43GAT), .B(G190GAT), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n411), .B(G134GAT), .ZN(n439) );
  XNOR2_X1 U479 ( .A(n439), .B(n412), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U481 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n566) );
  NAND2_X1 U485 ( .A1(n423), .A2(n566), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n424), .B(KEYINPUT47), .ZN(n430) );
  XNOR2_X1 U487 ( .A(KEYINPUT77), .B(n566), .ZN(n551) );
  INV_X1 U488 ( .A(n551), .ZN(n495) );
  XNOR2_X1 U489 ( .A(KEYINPUT36), .B(n495), .ZN(n589) );
  INV_X1 U490 ( .A(n570), .ZN(n586) );
  NOR2_X1 U491 ( .A1(n589), .A2(n586), .ZN(n425) );
  XNOR2_X1 U492 ( .A(KEYINPUT45), .B(n425), .ZN(n427) );
  NAND2_X1 U493 ( .A1(n427), .A2(n426), .ZN(n428) );
  NOR2_X1 U494 ( .A1(n428), .A2(n568), .ZN(n429) );
  NOR2_X1 U495 ( .A1(n430), .A2(n429), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n536) );
  AND2_X1 U497 ( .A1(n528), .A2(n536), .ZN(n435) );
  INV_X1 U498 ( .A(KEYINPUT120), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n574) );
  OR2_X1 U500 ( .A1(n292), .A2(n574), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n436), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT64), .Z(n442) );
  XOR2_X1 U503 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n438) );
  XNOR2_X1 U504 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n437) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n448) );
  XOR2_X1 U508 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U511 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n540) );
  NAND2_X1 U514 ( .A1(n453), .A2(n540), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n571), .A2(n558), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  NAND2_X1 U520 ( .A1(n568), .A2(n426), .ZN(n500) );
  XOR2_X1 U521 ( .A(n540), .B(KEYINPUT87), .Z(n462) );
  NAND2_X1 U522 ( .A1(n575), .A2(n468), .ZN(n537) );
  NOR2_X1 U523 ( .A1(n537), .A2(n542), .ZN(n460) );
  XNOR2_X1 U524 ( .A(KEYINPUT95), .B(n460), .ZN(n461) );
  NOR2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n477) );
  NAND2_X1 U526 ( .A1(n528), .A2(n540), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n463), .A2(n466), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n464), .B(KEYINPUT97), .ZN(n465) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n465), .Z(n471) );
  NOR2_X1 U530 ( .A1(n540), .A2(n466), .ZN(n467) );
  XNOR2_X1 U531 ( .A(KEYINPUT26), .B(n467), .ZN(n576) );
  AND2_X1 U532 ( .A1(n576), .A2(n468), .ZN(n469) );
  XNOR2_X1 U533 ( .A(KEYINPUT96), .B(n469), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n472), .B(KEYINPUT98), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n499) );
  NOR2_X1 U537 ( .A1(n499), .A2(n570), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n589), .A2(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(n481), .ZN(n526) );
  NOR2_X1 U540 ( .A1(n500), .A2(n526), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT38), .ZN(n511) );
  NAND2_X1 U542 ( .A1(n511), .A2(n540), .ZN(n484) );
  NAND2_X1 U543 ( .A1(n575), .A2(n511), .ZN(n488) );
  XOR2_X1 U544 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  AND2_X1 U547 ( .A1(n571), .A2(n551), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n490) );
  INV_X1 U549 ( .A(G190GAT), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n494) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n503) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n497) );
  NAND2_X1 U554 ( .A1(n570), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  OR2_X1 U556 ( .A1(n499), .A2(n498), .ZN(n513) );
  NOR2_X1 U557 ( .A1(n500), .A2(n513), .ZN(n501) );
  XNOR2_X1 U558 ( .A(KEYINPUT100), .B(n501), .ZN(n507) );
  NAND2_X1 U559 ( .A1(n575), .A2(n507), .ZN(n502) );
  XNOR2_X1 U560 ( .A(n503), .B(n502), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n507), .A2(n528), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n504), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT35), .Z(n506) );
  NAND2_X1 U564 ( .A1(n540), .A2(n507), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  XOR2_X1 U566 ( .A(G22GAT), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U567 ( .A1(n507), .A2(n542), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  NAND2_X1 U569 ( .A1(n511), .A2(n528), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n542), .ZN(n512) );
  XNOR2_X1 U572 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  INV_X1 U574 ( .A(n568), .ZN(n578) );
  NAND2_X1 U575 ( .A1(n578), .A2(n558), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n513), .A2(n525), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT106), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n575), .A2(n521), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  XOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT107), .Z(n518) );
  NAND2_X1 U581 ( .A1(n528), .A2(n521), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n540), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n520), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n542), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n575), .A2(n532), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n540), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT110), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n534) );
  NAND2_X1 U599 ( .A1(n532), .A2(n542), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  INV_X1 U602 ( .A(n536), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT114), .B(n539), .ZN(n556) );
  NAND2_X1 U605 ( .A1(n540), .A2(n556), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n568), .A2(n552), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U610 ( .A1(n552), .A2(n558), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT115), .Z(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U615 ( .A1(n552), .A2(n570), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(n555), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n576), .A2(n556), .ZN(n565) );
  NOR2_X1 U623 ( .A1(n578), .A2(n565), .ZN(n557) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n557), .Z(G1344GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n565), .A2(n559), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n561) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n586), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n571), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n578), .A2(n588), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n588), .A2(n426), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

