//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  OR2_X1    g006(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n218), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n210), .A2(new_n215), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT24), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n223), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(KEYINPUT24), .A3(new_n222), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT25), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n223), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n224), .ZN(new_n235));
  AND4_X1   g034(.A1(KEYINPUT25), .A2(new_n234), .A3(new_n235), .A4(new_n232), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n220), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G113gat), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g040(.A1(G113gat), .A2(G120gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n232), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n243), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n245), .B1(new_n243), .B2(KEYINPUT65), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n258), .A3(new_n220), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n205), .B1(new_n250), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G43gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G71gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G99gat), .ZN(new_n265));
  INV_X1    g064(.A(G71gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n263), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G99gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n205), .A3(new_n259), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n250), .A2(new_n274), .A3(new_n259), .A4(new_n205), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT33), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n265), .B2(new_n269), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(new_n281), .B(new_n286), .C1(new_n273), .C2(new_n275), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n262), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT34), .B1(new_n261), .B2(KEYINPUT68), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI211_X1 g090(.A(KEYINPUT69), .B(KEYINPUT34), .C1(new_n261), .C2(KEYINPUT68), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n286), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n262), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n278), .B1(new_n273), .B2(new_n275), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n295), .B(new_n296), .C1(new_n297), .C2(new_n271), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n288), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n293), .B1(new_n288), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n202), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n288), .A2(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(new_n293), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n293), .A3(new_n298), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT36), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n237), .A2(KEYINPUT71), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n255), .A2(new_n308), .A3(new_n220), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n307), .A2(G226gat), .A3(new_n309), .A4(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n237), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  INV_X1    g117(.A(G218gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n315), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n314), .B1(new_n255), .B2(new_n220), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n311), .A3(new_n309), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n313), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(new_n325), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  INV_X1    g130(.A(G64gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G92gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n326), .B(new_n335), .C1(new_n329), .C2(new_n325), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(G85gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(G155gat), .B2(G162gat), .ZN(new_n348));
  INV_X1    g147(.A(G148gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G141gat), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n348), .A2(KEYINPUT72), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n356));
  OR2_X1    g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n354), .A2(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n352), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n353), .A2(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n354), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n355), .A2(KEYINPUT72), .A3(KEYINPUT2), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n367), .A2(new_n361), .A3(new_n359), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n371), .A3(new_n258), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n373), .B(new_n375), .C1(new_n249), .C2(new_n363), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n249), .A2(new_n373), .A3(new_n363), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n258), .A2(new_n370), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n249), .A2(new_n363), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n383), .B2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(KEYINPUT73), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n249), .A2(new_n363), .A3(new_n387), .A4(new_n373), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT4), .B1(new_n258), .B2(new_n370), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n372), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n342), .B(new_n346), .C1(new_n385), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n385), .A2(new_n392), .ZN(new_n395));
  INV_X1    g194(.A(new_n346), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n385), .A2(new_n392), .A3(new_n346), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n342), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n339), .A2(new_n341), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n321), .A2(new_n323), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n322), .B1(new_n320), .B2(new_n316), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n311), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n364), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT75), .B1(new_n324), .B2(new_n311), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n370), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n365), .A2(new_n311), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n325), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n324), .B1(new_n365), .B2(new_n311), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n363), .B1(new_n405), .B2(new_n364), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n402), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT76), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n402), .A3(new_n417), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT74), .B(KEYINPUT31), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G78gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(G106gat), .Z(new_n425));
  NAND4_X1  g224(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n418), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n426), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n301), .A2(new_n306), .B1(new_n401), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n374), .B1(new_n390), .B2(new_n372), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n396), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n383), .A2(new_n375), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n372), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n389), .A2(new_n388), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n386), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT39), .B(new_n438), .C1(new_n441), .C2(new_n374), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n442), .A3(KEYINPUT40), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n397), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT40), .B1(new_n436), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(KEYINPUT77), .A3(new_n341), .A4(new_n339), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n339), .A2(new_n341), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n390), .A2(new_n372), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n435), .A3(new_n375), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n346), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n397), .A3(new_n443), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n448), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n330), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT37), .B(new_n326), .C1(new_n329), .C2(new_n325), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n335), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n398), .A2(new_n342), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n346), .B1(new_n385), .B2(new_n392), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n393), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n329), .A2(new_n325), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n310), .A2(new_n315), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(KEYINPUT37), .C1(new_n325), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n459), .A3(new_n470), .A4(new_n335), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n462), .A2(new_n466), .A3(new_n337), .A4(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n447), .A2(new_n457), .A3(new_n472), .A4(new_n431), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n299), .A2(new_n300), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n400), .A4(new_n431), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n304), .A2(new_n400), .A3(new_n431), .A4(new_n305), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n433), .A2(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT14), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT78), .B(G29gat), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G36gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT79), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT79), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(G36gat), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT15), .Z(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n491));
  INV_X1    g290(.A(new_n481), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n483), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  XOR2_X1   g295(.A(G15gat), .B(G22gat), .Z(new_n497));
  INV_X1    g296(.A(G1gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(G1gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT80), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G8gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n495), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n503), .B(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT81), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT17), .B(new_n493), .C1(new_n487), .C2(new_n489), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT82), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT82), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n510), .A2(new_n514), .A3(new_n519), .A4(new_n515), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n517), .A2(KEYINPUT84), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT11), .B(G169gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G197gat), .ZN(new_n523));
  XOR2_X1   g322(.A(G113gat), .B(G141gat), .Z(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  XOR2_X1   g324(.A(new_n525), .B(KEYINPUT12), .Z(new_n526));
  AND2_X1   g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n505), .A2(new_n509), .B1(new_n508), .B2(new_n506), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n515), .B(KEYINPUT83), .Z(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT13), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n516), .A2(new_n518), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n532), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n533), .ZN(new_n538));
  INV_X1    g337(.A(new_n526), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n479), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  AND3_X1   g343(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(KEYINPUT8), .A2(new_n546), .B1(new_n547), .B2(new_n334), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n547), .B2(new_n334), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n545), .B1(new_n495), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n512), .A2(new_n513), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n554), .ZN(new_n560));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561));
  AOI21_X1  g360(.A(new_n544), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n558), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n554), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n567), .A2(new_n568), .A3(new_n561), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  OAI22_X1  g369(.A1(new_n562), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n568), .ZN(new_n572));
  INV_X1    g371(.A(new_n561), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n560), .A2(new_n561), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n544), .A3(new_n575), .A4(new_n565), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G57gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G64gat), .ZN(new_n585));
  XOR2_X1   g384(.A(G71gat), .B(G78gat), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT86), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(new_n266), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n585), .A2(new_n587), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n586), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT20), .Z(new_n601));
  OAI21_X1  g400(.A(new_n508), .B1(new_n599), .B2(new_n598), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n602), .A2(G183gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(G183gat), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT88), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT89), .B(G211gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n605), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n582), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n581), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n578), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n621), .A3(new_n597), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n554), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n554), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT94), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(KEYINPUT95), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G176gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G204gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n598), .A2(new_n554), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT93), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n623), .A2(new_n625), .A3(KEYINPUT10), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n629), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(KEYINPUT95), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n634), .B1(new_n643), .B2(new_n630), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n619), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n543), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n466), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n498), .ZN(G1324gat));
  OAI21_X1  g449(.A(G8gat), .B1(new_n647), .B2(new_n449), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  INV_X1    g452(.A(new_n449), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT96), .B(G8gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  MUX2_X1   g456(.A(KEYINPUT42), .B(new_n652), .S(new_n657), .Z(G1325gat));
  NAND2_X1  g457(.A1(new_n301), .A2(new_n306), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(G15gat), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n474), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(G15gat), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT97), .Z(G1326gat));
  NOR2_X1   g464(.A1(new_n647), .A2(new_n431), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n666), .B(new_n668), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n578), .A2(new_n618), .A3(new_n645), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n543), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(new_n648), .A3(new_n482), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  OAI21_X1  g475(.A(KEYINPUT44), .B1(new_n479), .B2(new_n578), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n401), .A2(new_n432), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n473), .A2(new_n659), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n476), .A2(new_n478), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n577), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n618), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n645), .B(KEYINPUT100), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n684), .A2(new_n541), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n482), .B1(new_n687), .B2(new_n648), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n676), .A2(new_n688), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n687), .A2(new_n690), .A3(new_n449), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n687), .B2(new_n449), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(G36gat), .A3(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n674), .A2(G36gat), .A3(new_n449), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1329gat));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n674), .B2(new_n662), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n687), .A2(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n659), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g500(.A(new_n686), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n677), .B2(new_n683), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n541), .A3(new_n432), .A4(new_n685), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT102), .B1(new_n704), .B2(G50gat), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n674), .A2(G50gat), .A3(new_n431), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n704), .B2(G50gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n707), .B(new_n709), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n619), .A2(new_n686), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n681), .A2(new_n542), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n681), .A2(KEYINPUT103), .A3(new_n542), .A4(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n648), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT104), .B(G57gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1332gat));
  AND2_X1   g518(.A1(new_n714), .A2(new_n715), .ZN(new_n720));
  NAND2_X1  g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n654), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT105), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(KEYINPUT105), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n724), .A2(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1333gat));
  NAND3_X1  g529(.A1(new_n720), .A2(KEYINPUT106), .A3(new_n474), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n716), .B2(new_n662), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n266), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n720), .A2(G71gat), .A3(new_n660), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT50), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n716), .A2(new_n431), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(G78gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1335gat));
  INV_X1    g542(.A(new_n645), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n541), .A2(new_n618), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n744), .B(new_n746), .C1(new_n677), .C2(new_n683), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n648), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n479), .A2(new_n750), .A3(new_n746), .A4(new_n578), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n578), .B1(new_n679), .B2(new_n680), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n752), .B2(new_n745), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n744), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n547), .A3(new_n466), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n749), .A2(new_n756), .ZN(G1336gat));
  NOR3_X1   g556(.A1(new_n686), .A2(G92gat), .A3(new_n449), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n751), .B2(new_n753), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT109), .B(new_n758), .C1(new_n751), .C2(new_n753), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n684), .A2(new_n654), .A3(new_n645), .A4(new_n745), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(new_n764), .B2(G92gat), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(G92gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n681), .A2(new_n577), .A3(new_n745), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n750), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(new_n758), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n767), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT110), .B1(new_n766), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n774), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n763), .A2(new_n765), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n748), .B2(new_n659), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n755), .A2(new_n268), .A3(new_n474), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n748), .B2(new_n431), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n686), .A2(G106gat), .A3(new_n431), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n785), .C1(new_n754), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n786), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n790), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n792), .B2(new_n785), .ZN(G1339gat));
  INV_X1    g592(.A(new_n642), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n626), .A2(new_n636), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT93), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n637), .B(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n797), .A3(new_n628), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(new_n640), .A3(KEYINPUT54), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n800), .B(new_n629), .C1(new_n638), .C2(new_n639), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n634), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n804), .A3(new_n634), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n799), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n794), .B1(new_n806), .B2(KEYINPUT55), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(new_n805), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n804), .B1(new_n801), .B2(new_n634), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n799), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n541), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n510), .A2(new_n514), .ZN(new_n814));
  INV_X1    g613(.A(new_n515), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n814), .A2(new_n815), .B1(new_n528), .B2(new_n531), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n816), .B2(new_n525), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  INV_X1    g617(.A(new_n525), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n528), .A2(new_n531), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n515), .B1(new_n510), .B2(new_n514), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n527), .B2(new_n535), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n577), .B1(new_n824), .B2(new_n645), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n813), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n824), .A3(new_n812), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n577), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n685), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n646), .A2(new_n542), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n662), .A2(new_n432), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n654), .A2(new_n648), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n541), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g637(.A(new_n239), .B1(new_n836), .B2(new_n702), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n645), .A2(new_n239), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT114), .Z(new_n841));
  AOI21_X1  g640(.A(new_n839), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n842), .B(new_n843), .ZN(G1341gat));
  NAND3_X1  g643(.A1(new_n836), .A2(G127gat), .A3(new_n618), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  AOI21_X1  g647(.A(G127gat), .B1(new_n836), .B2(new_n618), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1342gat));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n833), .A2(new_n578), .A3(new_n835), .ZN(new_n852));
  INV_X1    g651(.A(G134gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n618), .B1(new_n813), .B2(new_n825), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n855), .A2(new_n828), .B1(new_n646), .B2(new_n542), .ZN(new_n856));
  INV_X1    g655(.A(new_n832), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n577), .A3(new_n834), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT56), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n854), .A2(new_n860), .A3(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(G134gat), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n854), .C2(new_n860), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(G1343gat));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n856), .B2(new_n431), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n831), .A2(new_n869), .A3(new_n432), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n660), .A2(new_n835), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n870), .A3(new_n541), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n542), .A2(G141gat), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n432), .A2(new_n831), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT119), .B1(new_n872), .B2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n873), .B2(new_n876), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT120), .B(new_n875), .C1(new_n872), .C2(G141gat), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n884), .A2(new_n885), .B1(KEYINPUT58), .B2(new_n879), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(G1344gat));
  AND3_X1   g686(.A1(new_n831), .A2(new_n432), .A3(new_n871), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n349), .A3(new_n645), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n870), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n645), .A3(new_n871), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(G148gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  AOI21_X1  g695(.A(G155gat), .B1(new_n888), .B2(new_n618), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n890), .A2(new_n660), .A3(new_n835), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n618), .A2(G155gat), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT121), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n888), .B2(new_n577), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n898), .A2(new_n577), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n449), .A2(new_n466), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n474), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n432), .B1(new_n906), .B2(KEYINPUT122), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n831), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n542), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n858), .A2(new_n905), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n226), .A3(new_n541), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1348gat));
  NOR3_X1   g713(.A1(new_n910), .A2(new_n227), .A3(new_n686), .ZN(new_n915));
  AOI21_X1  g714(.A(G176gat), .B1(new_n912), .B2(new_n645), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  AOI21_X1  g716(.A(new_n230), .B1(new_n909), .B2(new_n618), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n618), .A2(new_n206), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g720(.A(new_n207), .B1(new_n909), .B2(new_n577), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n207), .A3(new_n577), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1351gat));
  OR2_X1    g725(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n659), .A2(new_n905), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n542), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n659), .A2(new_n654), .A3(new_n432), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n466), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n831), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(G197gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n931), .B1(new_n542), .B2(new_n938), .ZN(G1352gat));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(G204gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n930), .B2(new_n686), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n937), .A2(new_n744), .A3(new_n940), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n936), .A2(new_n318), .A3(new_n618), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n891), .A2(new_n618), .A3(new_n928), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  NAND2_X1  g748(.A1(new_n577), .A2(G218gat), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n319), .B1(new_n937), .B2(new_n578), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(G1355gat));
endmodule


