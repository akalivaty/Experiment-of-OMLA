//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923;
  INV_X1    g000(.A(G148gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT75), .B1(new_n202), .B2(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n206), .C1(new_n205), .C2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n202), .A2(G141gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n205), .A2(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n209), .A2(new_n208), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221));
  XNOR2_X1  g020(.A(G197gat), .B(G204gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT22), .ZN(new_n223));
  INV_X1    g022(.A(G211gat), .ZN(new_n224));
  INV_X1    g023(.A(G218gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n221), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n217), .A3(new_n221), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n230), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n220), .A2(new_n232), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n229), .B2(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n218), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n229), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(G22gat), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G22gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(new_n242), .C1(new_n235), .C2(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(KEYINPUT78), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT31), .ZN(new_n249));
  INV_X1    g048(.A(G50gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n251), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n254), .A4(new_n246), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n244), .A2(new_n254), .A3(new_n246), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(new_n258), .A3(KEYINPUT80), .A4(new_n255), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g066(.A1(G113gat), .A2(G120gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT67), .B1(new_n269), .B2(KEYINPUT68), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g072(.A(new_n271), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(KEYINPUT67), .C1(new_n269), .C2(KEYINPUT68), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(G183gat), .A3(G190gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G183gat), .B(G190gat), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT65), .B(new_n278), .C1(new_n279), .C2(new_n277), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT23), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n280), .B(new_n281), .C1(new_n282), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n278), .ZN(new_n291));
  INV_X1    g090(.A(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G190gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n291), .B1(new_n296), .B2(KEYINPUT24), .ZN(new_n297));
  INV_X1    g096(.A(new_n289), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n297), .B(new_n298), .C1(KEYINPUT65), .C2(KEYINPUT25), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(KEYINPUT27), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n303), .A3(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n283), .A3(new_n284), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n288), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n301), .A2(new_n303), .A3(new_n311), .A4(new_n294), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n305), .A2(new_n306), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n309), .A2(new_n288), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n316), .A2(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n317), .A2(KEYINPUT66), .A3(new_n305), .A4(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n276), .B1(new_n300), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n321), .B(KEYINPUT64), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n290), .A2(new_n299), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n315), .A4(new_n318), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT33), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(KEYINPUT69), .A3(new_n327), .ZN(new_n331));
  XNOR2_X1  g130(.A(G15gat), .B(G43gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n326), .B2(KEYINPUT32), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n326), .B(KEYINPUT32), .C1(new_n327), .C2(new_n334), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n325), .ZN(new_n339));
  INV_X1    g138(.A(new_n322), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT34), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT70), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n344), .A3(KEYINPUT34), .ZN(new_n345));
  AOI211_X1 g144(.A(KEYINPUT34), .B(new_n322), .C1(new_n320), .C2(new_n325), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n342), .B2(KEYINPUT70), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n336), .A2(new_n350), .A3(new_n337), .A4(new_n345), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n263), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n323), .A2(new_n313), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n315), .A3(new_n318), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n231), .A2(new_n355), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n353), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n229), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n360));
  OAI22_X1  g159(.A1(new_n353), .A2(new_n360), .B1(new_n356), .B2(new_n354), .ZN(new_n361));
  INV_X1    g160(.A(new_n229), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G64gat), .ZN(new_n365));
  INV_X1    g164(.A(G92gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n359), .A2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n352), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n324), .A3(new_n233), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n218), .B(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n276), .ZN(new_n384));
  INV_X1    g183(.A(new_n218), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n276), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n324), .A2(new_n218), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n381), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n383), .A2(new_n387), .A3(new_n276), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n390), .A3(new_n382), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(G57gat), .ZN(new_n403));
  INV_X1    g202(.A(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n378), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n406), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n378), .C1(new_n400), .C2(new_n406), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT35), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n351), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n338), .A2(new_n418), .A3(new_n348), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n409), .A2(new_n378), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n400), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n405), .B(KEYINPUT82), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT84), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n407), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n376), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n263), .A2(new_n420), .A3(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n377), .A2(new_n416), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n381), .B1(new_n398), .B2(new_n380), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n392), .A2(new_n393), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n435), .B2(KEYINPUT83), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(KEYINPUT83), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT40), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n426), .A3(new_n376), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n372), .B1(new_n371), .B2(KEYINPUT37), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n359), .B2(new_n363), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT38), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n358), .B2(new_n362), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n361), .A2(new_n229), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT38), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n369), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n263), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n376), .B1(new_n412), .B2(new_n413), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n263), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n417), .A2(new_n454), .A3(new_n419), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n349), .A2(KEYINPUT36), .A3(new_n351), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n349), .A2(KEYINPUT71), .A3(new_n351), .A4(KEYINPUT36), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n455), .A2(KEYINPUT73), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n417), .A2(new_n461), .A3(new_n454), .A4(new_n419), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n453), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n451), .B1(new_n463), .B2(KEYINPUT81), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n453), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT81), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n431), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n473));
  INV_X1    g272(.A(G1gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT89), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G1gat), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n471), .A2(G1gat), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n481), .A2(G8gat), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(G8gat), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G78gat), .ZN(new_n486));
  INV_X1    g285(.A(G57gat), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n487), .A2(G64gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(G64gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n490), .B2(KEYINPUT9), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n486), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494));
  INV_X1    g293(.A(G71gat), .ZN(new_n495));
  INV_X1    g294(.A(G78gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n489), .A2(KEYINPUT92), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(KEYINPUT92), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n488), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n493), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT94), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n493), .A2(new_n503), .A3(new_n497), .A4(new_n500), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n485), .B1(KEYINPUT21), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(new_n292), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n508));
  NAND2_X1  g307(.A1(G231gat), .A2(G233gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n507), .B(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n505), .A2(KEYINPUT21), .ZN(new_n512));
  XNOR2_X1  g311(.A(G127gat), .B(G155gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n224), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n511), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT97), .ZN(new_n518));
  AND2_X1   g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT41), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n518), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT86), .B(G29gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT87), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  INV_X1    g325(.A(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT14), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G43gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G50gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n535), .A2(G50gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n538), .B1(new_n542), .B2(new_n536), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n542), .B2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n539), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n540), .A2(new_n531), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n541), .A2(KEYINPUT17), .A3(new_n547), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT95), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n404), .B2(new_n366), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n554), .A2(new_n559), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n563), .A2(new_n548), .B1(KEYINPUT41), .B2(new_n519), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n565), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n522), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n566), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n521), .A3(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  OR3_X1    g375(.A1(new_n516), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT98), .B1(new_n516), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT11), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n283), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G197gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT12), .ZN(new_n584));
  INV_X1    g383(.A(new_n485), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n550), .A3(new_n551), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n586), .A2(new_n587), .B1(new_n485), .B2(new_n548), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n485), .B(new_n548), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n590), .B(KEYINPUT13), .Z(new_n594));
  AOI22_X1  g393(.A1(new_n591), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT18), .A4(new_n590), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n584), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n594), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n584), .A3(new_n596), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n560), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT99), .B1(new_n554), .B2(new_n559), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n505), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n563), .B2(new_n505), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT101), .Z(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT100), .B(KEYINPUT10), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n607), .B(new_n613), .C1(new_n563), .C2(new_n505), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n563), .A2(KEYINPUT10), .A3(new_n505), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G176gat), .ZN(new_n619));
  INV_X1    g418(.A(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n611), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n579), .A2(new_n603), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n470), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n414), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G8gat), .Z(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n376), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n376), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G8gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n628), .A2(new_n639), .A3(new_n420), .ZN(new_n640));
  INV_X1    g439(.A(new_n467), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n642), .B2(new_n639), .ZN(G1326gat));
  INV_X1    g442(.A(new_n263), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT102), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n645), .B(new_n647), .ZN(G1327gat));
  INV_X1    g447(.A(new_n516), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n603), .A2(new_n649), .A3(new_n626), .ZN(new_n650));
  INV_X1    g449(.A(new_n576), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n463), .A2(new_n451), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n431), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n470), .B2(new_n576), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(KEYINPUT103), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n658), .B(new_n654), .C1(new_n470), .C2(new_n576), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n650), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(new_n650), .C1(new_n657), .C2(new_n659), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n414), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n661), .A2(KEYINPUT105), .A3(new_n414), .A4(new_n663), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n523), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n470), .A2(new_n576), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n650), .ZN(new_n670));
  INV_X1    g469(.A(new_n414), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n670), .A2(new_n671), .A3(new_n523), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT45), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(G1328gat));
  INV_X1    g473(.A(new_n376), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n670), .A2(G36gat), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT46), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n661), .A2(new_n376), .A3(new_n663), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n527), .ZN(G1329gat));
  OAI21_X1  g478(.A(G43gat), .B1(new_n660), .B2(new_n467), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n669), .A2(new_n535), .A3(new_n420), .A4(new_n650), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(KEYINPUT47), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n641), .A3(new_n663), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(G43gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n682), .B1(new_n685), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g485(.A1(new_n670), .A2(G50gat), .A3(new_n263), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n660), .B2(new_n263), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G50gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n660), .A2(new_n690), .A3(new_n263), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n661), .A2(new_n644), .A3(new_n663), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n687), .B1(new_n695), .B2(G50gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g496(.A(new_n626), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n579), .A2(new_n602), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n431), .A2(new_n652), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n671), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n487), .ZN(G1332gat));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n675), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  AND2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n701), .B2(new_n467), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n420), .A2(new_n495), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g511(.A1(new_n701), .A2(new_n263), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n496), .ZN(G1335gat));
  OR2_X1    g513(.A1(new_n657), .A2(new_n659), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n649), .A2(new_n602), .A3(new_n698), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717), .B2(new_n671), .ZN(new_n718));
  INV_X1    g517(.A(new_n653), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n603), .B(new_n516), .C1(new_n653), .C2(KEYINPUT107), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT51), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n721), .B2(new_n722), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n698), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n404), .A3(new_n414), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n718), .A2(new_n728), .ZN(G1336gat));
  NOR2_X1   g528(.A1(new_n675), .A2(G92gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n376), .B(new_n716), .C1(new_n657), .C2(new_n659), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G92gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n733), .A2(new_n736), .A3(G92gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n733), .B2(G92gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n626), .A2(new_n730), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n723), .B1(KEYINPUT109), .B2(KEYINPUT51), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n721), .B2(new_n722), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n735), .B1(new_n744), .B2(new_n732), .ZN(G1337gat));
  INV_X1    g544(.A(G99gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n717), .A2(new_n746), .A3(new_n467), .ZN(new_n747));
  AOI21_X1  g546(.A(G99gat), .B1(new_n727), .B2(new_n420), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1338gat));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n715), .A2(new_n644), .A3(new_n716), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n740), .A2(new_n742), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n698), .A2(G106gat), .A3(new_n263), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT110), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n751), .A2(G106gat), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n751), .A2(G106gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n724), .A2(new_n726), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n753), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n750), .A2(new_n755), .B1(new_n756), .B2(new_n759), .ZN(G1339gat));
  NAND4_X1  g559(.A1(new_n577), .A2(new_n603), .A3(new_n578), .A4(new_n698), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n590), .B1(new_n588), .B2(new_n589), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n593), .A2(new_n594), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n583), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n576), .A2(new_n601), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n614), .A2(new_n610), .A3(new_n615), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n617), .A2(KEYINPUT54), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n616), .A2(new_n768), .A3(new_n609), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(new_n624), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n624), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT55), .B(new_n767), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n765), .A2(new_n775), .A3(new_n622), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n776), .A2(new_n622), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n775), .A4(new_n765), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n626), .A2(new_n601), .A3(new_n764), .ZN(new_n782));
  INV_X1    g581(.A(new_n601), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n776), .B(new_n622), .C1(new_n783), .C2(new_n597), .ZN(new_n784));
  INV_X1    g583(.A(new_n775), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n778), .A2(new_n781), .B1(new_n786), .B2(new_n651), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n761), .B1(new_n787), .B2(new_n649), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(new_n263), .A3(new_n420), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n671), .A2(new_n376), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(new_n264), .A3(new_n603), .ZN(new_n792));
  INV_X1    g591(.A(new_n788), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n671), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n377), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n602), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n792), .B1(new_n797), .B2(new_n264), .ZN(G1340gat));
  OAI21_X1  g597(.A(G120gat), .B1(new_n791), .B2(new_n698), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n265), .A3(new_n626), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n791), .A2(new_n803), .A3(new_n516), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n649), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n805), .A2(KEYINPUT115), .ZN(new_n806));
  AOI21_X1  g605(.A(G127gat), .B1(new_n805), .B2(KEYINPUT115), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(G1342gat));
  NOR2_X1   g607(.A1(new_n651), .A2(G134gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n377), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n789), .A2(new_n576), .A3(new_n790), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(G134gat), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n810), .B2(KEYINPUT56), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n810), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n813), .B(KEYINPUT117), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1343gat));
  NOR3_X1   g619(.A1(new_n641), .A2(new_n263), .A3(new_n376), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n794), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n205), .A3(new_n602), .ZN(new_n824));
  XOR2_X1   g623(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n825));
  NAND2_X1  g624(.A1(new_n773), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n779), .A2(new_n602), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n576), .B1(new_n827), .B2(new_n782), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT119), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n828), .A2(KEYINPUT119), .B1(new_n778), .B2(new_n781), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n649), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n761), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n644), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n788), .A2(new_n835), .A3(new_n644), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n467), .A2(new_n790), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n603), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n824), .B1(new_n841), .B2(new_n205), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT58), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n202), .A2(KEYINPUT59), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n840), .B2(new_n698), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n835), .B1(new_n788), .B2(new_n644), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n644), .A2(new_n835), .ZN(new_n849));
  INV_X1    g648(.A(new_n777), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n516), .B1(new_n828), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n761), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n788), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n644), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n626), .A3(new_n838), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n846), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n858), .B(new_n846), .C1(new_n855), .C2(G148gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n845), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n823), .A2(new_n202), .A3(new_n626), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1345gat));
  OAI21_X1  g661(.A(G155gat), .B1(new_n840), .B2(new_n516), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n516), .A2(G155gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n822), .B2(new_n864), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n840), .B2(new_n651), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n651), .A2(G162gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n822), .B2(new_n867), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n414), .A2(new_n675), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n789), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n283), .A3(new_n603), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n793), .A2(new_n414), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n352), .A2(new_n675), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n602), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(new_n283), .ZN(G1348gat));
  OAI21_X1  g676(.A(G176gat), .B1(new_n870), .B2(new_n698), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n626), .A2(new_n284), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n874), .B2(new_n879), .ZN(G1349gat));
  OAI21_X1  g679(.A(G183gat), .B1(new_n870), .B2(new_n516), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n649), .A2(new_n301), .A3(new_n303), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g683(.A1(new_n875), .A2(new_n294), .A3(new_n576), .ZN(new_n885));
  OAI21_X1  g684(.A(G190gat), .B1(new_n870), .B2(new_n651), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT61), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(KEYINPUT61), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT123), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n885), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n641), .A2(new_n263), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n376), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT124), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n872), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(G197gat), .A3(new_n603), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n467), .A2(new_n869), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT126), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n853), .A2(new_n854), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G197gat), .B1(new_n903), .B2(new_n603), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n853), .A2(new_n626), .A3(new_n854), .ZN(new_n906));
  OAI21_X1  g705(.A(G204gat), .B1(new_n906), .B2(new_n901), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n698), .A2(G204gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n897), .B2(new_n909), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n897), .A2(KEYINPUT62), .A3(new_n909), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(G1353gat));
  INV_X1    g711(.A(new_n897), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n224), .A3(new_n649), .ZN(new_n914));
  OAI21_X1  g713(.A(G211gat), .B1(new_n903), .B2(new_n516), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1354gat));
  AND2_X1   g718(.A1(new_n903), .A2(KEYINPUT127), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n576), .B1(new_n903), .B2(KEYINPUT127), .ZN(new_n921));
  OAI21_X1  g720(.A(G218gat), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n913), .A2(new_n225), .A3(new_n576), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1355gat));
endmodule


