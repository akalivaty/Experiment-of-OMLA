//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n215), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT64), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n245), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G77), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n204), .A2(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n212), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n246), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n252), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n254), .A2(new_n258), .A3(new_n259), .A4(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(G274), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G226), .A2(G1698), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n227), .B2(G1698), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(G33), .B2(G97), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n270), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(G238), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n266), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n269), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT72), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n276), .A2(new_n277), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n282), .A2(new_n285), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT13), .B1(new_n288), .B2(new_n275), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT14), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G169), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n287), .A2(new_n289), .A3(G179), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n290), .B2(G169), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n263), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(new_n263), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n290), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(new_n301), .B(KEYINPUT73), .Z(new_n302));
  INV_X1    g0102(.A(new_n260), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n261), .A2(G50), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n303), .A2(new_n304), .B1(G50), .B2(new_n255), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G50), .A2(G58), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n204), .B1(new_n306), .B2(new_n246), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT8), .B(G58), .ZN(new_n308));
  INV_X1    g0108(.A(G150), .ZN(new_n309));
  INV_X1    g0109(.A(new_n245), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n308), .A2(new_n249), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(KEYINPUT69), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(KEYINPUT69), .B2(new_n311), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n305), .B1(new_n313), .B2(new_n252), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT68), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n273), .A2(new_n323), .A3(G1698), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n315), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n273), .A2(new_n321), .ZN(new_n326));
  INV_X1    g0126(.A(G222), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(new_n248), .B2(new_n273), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n283), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n270), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G226), .B2(new_n284), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G179), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n314), .B(new_n333), .C1(new_n334), .C2(new_n332), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n313), .A2(new_n252), .ZN(new_n336));
  INV_X1    g0136(.A(new_n305), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n338), .A2(new_n339), .B1(new_n332), .B2(new_n299), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT10), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n332), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G190), .B1(new_n314), .B2(KEYINPUT9), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n341), .A4(new_n340), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n335), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n315), .A2(new_n321), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G1698), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n317), .A2(new_n350), .A3(new_n319), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n283), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n266), .A2(G232), .A3(new_n279), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n270), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n266), .B1(new_n353), .B2(new_n354), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n270), .A2(new_n357), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n334), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n360), .B2(new_n364), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n308), .B1(new_n203), .B2(G20), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n260), .B1(new_n256), .B2(new_n308), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n252), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n246), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n245), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n320), .A2(new_n204), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n246), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n320), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT7), .A2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n377), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n371), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT75), .B1(new_n318), .B2(G33), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n316), .A3(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(new_n319), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n273), .B2(G20), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n246), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n387), .B1(new_n396), .B2(new_n377), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n370), .B1(new_n386), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT18), .B1(new_n367), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n377), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT74), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT74), .B1(new_n317), .B2(new_n319), .ZN(new_n402));
  INV_X1    g0202(.A(new_n383), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(G20), .B1(new_n317), .B2(new_n319), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n405), .B2(new_n392), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n400), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n252), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n394), .A2(new_n395), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT16), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n369), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(G169), .B1(new_n356), .B2(new_n358), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n362), .A2(new_n363), .A3(G179), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT76), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n360), .A2(new_n364), .A3(new_n361), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G200), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n356), .B2(new_n358), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT77), .B(G190), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n362), .A2(new_n363), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n369), .C1(new_n408), .C2(new_n411), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n399), .A2(new_n419), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n322), .A2(new_n324), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G238), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n326), .A2(new_n227), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT70), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G107), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n273), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n266), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G244), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n270), .B1(new_n280), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n359), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n334), .B1(new_n442), .B2(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n261), .A2(G77), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n303), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n248), .B2(new_n256), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n310), .A2(KEYINPUT71), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n310), .A2(KEYINPUT71), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n452), .A2(new_n308), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n455), .A2(new_n249), .B1(new_n204), .B2(new_n248), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n252), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n450), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n446), .A2(new_n447), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n445), .A2(G190), .ZN(new_n460));
  OAI21_X1  g0260(.A(G200), .B1(new_n442), .B2(new_n444), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n457), .A3(new_n450), .A4(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n349), .A2(new_n430), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n302), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n434), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT25), .B1(new_n256), .B2(new_n434), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n203), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n255), .A2(new_n469), .A3(new_n212), .A4(new_n251), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n467), .A2(new_n468), .B1(new_n434), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  INV_X1    g0274(.A(G250), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n326), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n283), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n268), .A2(G1), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n283), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G264), .ZN(new_n481));
  INV_X1    g0281(.A(G274), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n264), .B2(new_n265), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(new_n478), .A3(new_n479), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n420), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n476), .A2(new_n283), .B1(G264), .B2(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n299), .A3(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n438), .B2(new_n204), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT80), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n204), .A3(G33), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n434), .A3(G20), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(new_n434), .A3(KEYINPUT85), .A4(G20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n491), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n317), .A2(new_n319), .A3(new_n204), .A4(G87), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n273), .A2(KEYINPUT22), .A3(new_n204), .A4(G87), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n491), .A2(new_n503), .A3(new_n497), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT24), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT86), .B1(new_n515), .B2(new_n252), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n517), .B(new_n371), .C1(new_n511), .C2(new_n514), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n472), .B(new_n489), .C1(new_n516), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n510), .B1(new_n504), .B2(new_n509), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT24), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n252), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n252), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n471), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n485), .A2(new_n334), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(G179), .B2(new_n485), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT21), .ZN(new_n529));
  AND2_X1   g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n478), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n480), .A2(G270), .B1(new_n533), .B2(new_n483), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n317), .A2(new_n319), .A3(G264), .A4(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n317), .A2(new_n319), .A3(G257), .A4(new_n321), .ZN(new_n536));
  INV_X1    g0336(.A(G303), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n273), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n283), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n470), .A2(new_n492), .B1(new_n496), .B2(new_n255), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  AOI21_X1  g0343(.A(G20), .B1(G33), .B2(G283), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n316), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n252), .B1(new_n496), .B2(new_n204), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n493), .A2(new_n495), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n371), .B1(new_n552), .B2(G20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n545), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT83), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n557), .A3(KEYINPUT20), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n542), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n529), .B1(new_n541), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n542), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n549), .A2(new_n543), .A3(new_n550), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT20), .B1(new_n553), .B2(new_n557), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n334), .B1(new_n534), .B2(new_n539), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(KEYINPUT21), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n538), .A2(new_n283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n532), .A2(new_n266), .ZN(new_n568));
  INV_X1    g0368(.A(G270), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n484), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n422), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n534), .A2(new_n539), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n559), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n534), .A2(new_n539), .A3(G179), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n564), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n560), .A2(new_n566), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n317), .A2(new_n319), .A3(G244), .A4(new_n321), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n321), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G283), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n283), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n532), .A2(G257), .A3(new_n266), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n484), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G179), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n589), .A3(KEYINPUT79), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n585), .B2(new_n283), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n592), .A2(new_n593), .B1(new_n334), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G97), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n256), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n470), .B2(new_n597), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n597), .A2(new_n434), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G97), .A2(G107), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n434), .A2(KEYINPUT6), .A3(G97), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n245), .A2(G77), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n378), .A2(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n439), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT78), .B1(new_n611), .B2(new_n252), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n439), .B1(new_n394), .B2(new_n395), .ZN(new_n613));
  XNOR2_X1  g0413(.A(G97), .B(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n605), .B1(new_n614), .B2(new_n601), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n204), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT78), .B(new_n252), .C1(new_n613), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n600), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n596), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n252), .B1(new_n613), .B2(new_n616), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT78), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n599), .B1(new_n623), .B2(new_n617), .ZN(new_n624));
  INV_X1    g0424(.A(new_n588), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n586), .A2(new_n299), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G200), .B2(new_n594), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n494), .A2(G116), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n492), .A2(KEYINPUT80), .ZN(new_n630));
  OAI21_X1  g0430(.A(G33), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n278), .A2(new_n321), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n443), .A2(G1698), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n317), .A2(new_n632), .A3(new_n319), .A4(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n266), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n266), .A2(G274), .A3(new_n478), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n475), .B1(new_n203), .B2(G45), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n266), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n483), .A2(new_n478), .B1(new_n266), .B2(new_n637), .ZN(new_n641));
  NOR2_X1   g0441(.A1(G238), .A2(G1698), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n443), .B2(G1698), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n273), .B1(new_n496), .B2(G33), .ZN(new_n644));
  OAI211_X1 g0444(.A(G179), .B(new_n641), .C1(new_n644), .C2(new_n266), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n455), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n255), .ZN(new_n648));
  NOR2_X1   g0448(.A1(G87), .A2(G97), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n435), .A2(new_n437), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n204), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT19), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT81), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n317), .A2(new_n319), .A3(new_n204), .A4(G68), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n654), .A2(KEYINPUT81), .A3(new_n655), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n653), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n648), .B1(new_n661), .B2(new_n252), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n260), .A2(KEYINPUT82), .A3(new_n469), .A4(new_n647), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT82), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n470), .B2(new_n455), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G87), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n470), .A2(new_n668), .ZN(new_n669));
  AOI211_X1 g0469(.A(new_n648), .B(new_n669), .C1(new_n661), .C2(new_n252), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n420), .B1(new_n635), .B2(new_n639), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n299), .B(new_n641), .C1(new_n644), .C2(new_n266), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n646), .A2(new_n667), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n578), .A2(new_n620), .A3(new_n628), .A4(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n465), .A2(new_n528), .A3(new_n675), .ZN(G372));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n646), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n673), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n519), .A3(new_n620), .A4(new_n628), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n560), .A2(new_n577), .A3(new_n566), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n472), .B1(new_n516), .B2(new_n518), .ZN(new_n685));
  INV_X1    g0485(.A(new_n527), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n596), .A2(new_n619), .A3(new_n674), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n671), .A2(new_n672), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n661), .A2(new_n252), .ZN(new_n692));
  INV_X1    g0492(.A(new_n648), .ZN(new_n693));
  INV_X1    g0493(.A(new_n669), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n662), .A2(new_n666), .B1(new_n640), .B2(new_n645), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT87), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n619), .A3(new_n596), .A4(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n690), .B(new_n677), .C1(new_n700), .C2(KEYINPUT26), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n464), .B1(new_n688), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n344), .A2(new_n348), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n459), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT88), .A4(new_n458), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n300), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n296), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n427), .A2(new_n428), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n399), .A2(new_n419), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n703), .B1(new_n712), .B2(KEYINPUT89), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT89), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n335), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n702), .A2(new_n716), .ZN(G369));
  NAND3_X1  g0517(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT90), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT27), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT90), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n203), .A3(new_n204), .A4(G13), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT91), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n719), .A2(KEYINPUT91), .A3(new_n720), .A4(new_n722), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G213), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n719), .A2(new_n722), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(KEYINPUT27), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n727), .A2(G343), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n564), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n578), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n684), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n732), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  INV_X1    g0536(.A(new_n731), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n525), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n685), .A2(new_n686), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n528), .A2(new_n738), .B1(new_n739), .B2(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n685), .A2(new_n686), .A3(new_n737), .ZN(new_n742));
  INV_X1    g0542(.A(new_n528), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n734), .A2(new_n731), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(G399));
  INV_X1    g0546(.A(new_n207), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n650), .A2(G116), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(G1), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n210), .B2(new_n749), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n675), .A2(new_n528), .A3(new_n731), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n635), .A2(new_n639), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n487), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT92), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n756), .A2(new_n576), .A3(new_n594), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n594), .A2(new_n487), .A3(new_n755), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n761), .B2(new_n575), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n755), .A2(G179), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n595), .A2(new_n485), .A3(new_n540), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT31), .B1(new_n765), .B2(new_n731), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G330), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n737), .B1(new_n688), .B2(new_n701), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT93), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT29), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT93), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n776), .B(new_n737), .C1(new_n688), .C2(new_n701), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT26), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n596), .A2(new_n619), .A3(new_n779), .A4(new_n674), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n677), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(KEYINPUT26), .B2(new_n700), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n734), .B1(new_n525), .B2(new_n527), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n586), .A2(new_n589), .A3(KEYINPUT79), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT79), .B1(new_n586), .B2(new_n589), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G169), .B2(new_n594), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n624), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n623), .A2(new_n617), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n788), .A2(new_n627), .A3(new_n600), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n783), .A2(new_n790), .A3(new_n519), .A4(new_n682), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n731), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT29), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n772), .B1(new_n778), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n753), .B1(new_n794), .B2(G1), .ZN(G364));
  INV_X1    g0595(.A(G13), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G45), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT94), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n800), .A2(new_n748), .A3(new_n203), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT95), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n212), .B1(G20), .B2(new_n334), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G179), .A2(G200), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n204), .B1(new_n808), .B2(G190), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n597), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT98), .B1(new_n420), .B2(G179), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n420), .A2(KEYINPUT98), .A3(G179), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n204), .A2(new_n299), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n299), .A2(G20), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT97), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n817), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n273), .B1(new_n820), .B2(new_n668), .C1(new_n825), .C2(new_n434), .ZN(new_n826));
  NAND2_X1  g0626(.A1(G20), .A2(G179), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n420), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n422), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n813), .B(new_n826), .C1(G58), .C2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n823), .A2(G179), .A3(G200), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n833), .A2(KEYINPUT32), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n829), .A2(G190), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G50), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n828), .A2(new_n572), .A3(G200), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n837), .A2(new_n248), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT32), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n832), .B2(G159), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n835), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n828), .A2(new_n299), .A3(G200), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT99), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n831), .B(new_n843), .C1(new_n246), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n820), .B(KEYINPUT101), .Z(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G303), .ZN(new_n851));
  INV_X1    g0651(.A(new_n848), .ZN(new_n852));
  XNOR2_X1  g0652(.A(KEYINPUT33), .B(G317), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n830), .ZN(new_n855));
  INV_X1    g0655(.A(G322), .ZN(new_n856));
  INV_X1    g0656(.A(G326), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(new_n839), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  INV_X1    g0659(.A(G294), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n837), .A2(new_n859), .B1(new_n860), .B2(new_n812), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n320), .B1(new_n825), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G329), .B2(new_n832), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n851), .A2(new_n854), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n807), .B1(new_n849), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(G13), .A2(G33), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(G20), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(new_n806), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n401), .A2(new_n402), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n207), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n268), .B2(new_n211), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n240), .B2(new_n268), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n747), .A2(new_n320), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(G355), .B1(new_n492), .B2(new_n747), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n805), .B(new_n867), .C1(new_n871), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n870), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n735), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT102), .ZN(new_n882));
  INV_X1    g0682(.A(new_n805), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n736), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(G330), .B2(new_n735), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(G396));
  NAND4_X1  g0686(.A1(new_n705), .A2(new_n458), .A3(new_n706), .A4(new_n731), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n458), .A2(new_n731), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n462), .A2(new_n459), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n774), .A2(new_n777), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n737), .C1(new_n688), .C2(new_n701), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n772), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n803), .B2(new_n804), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n772), .A3(new_n893), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n806), .A2(new_n868), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n805), .B1(new_n248), .B2(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n860), .A2(new_n855), .B1(new_n837), .B2(new_n552), .ZN(new_n900));
  INV_X1    g0700(.A(new_n839), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n813), .B(new_n900), .C1(G303), .C2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n320), .B1(new_n833), .B2(new_n859), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(G87), .B2(new_n824), .ZN(new_n904));
  INV_X1    g0704(.A(new_n850), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n902), .B(new_n904), .C1(new_n434), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n848), .A2(new_n863), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n836), .A2(G159), .B1(new_n901), .B2(G137), .ZN(new_n909));
  INV_X1    g0709(.A(G143), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n909), .B1(new_n910), .B2(new_n855), .C1(new_n848), .C2(new_n309), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT34), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n872), .B1(new_n832), .B2(G132), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n824), .A2(G68), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(new_n372), .C2(new_n812), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n850), .B2(G50), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n908), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n899), .B1(new_n890), .B2(new_n869), .C1(new_n807), .C2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n897), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(G384));
  OR2_X1    g0720(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(G116), .A4(new_n213), .ZN(new_n923));
  XNOR2_X1  g0723(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(G77), .B1(new_n372), .B2(new_n246), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n927), .A2(new_n210), .B1(G50), .B2(new_n246), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n796), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT104), .ZN(new_n931));
  INV_X1    g0731(.A(new_n295), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n300), .A2(new_n932), .A3(new_n293), .A4(new_n292), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n263), .A2(new_n731), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(KEYINPUT105), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n296), .A2(new_n300), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n459), .A2(new_n731), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n893), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT38), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT37), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n727), .A2(new_n730), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n412), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n412), .A2(new_n417), .ZN(new_n950));
  AND4_X1   g0750(.A1(new_n945), .A2(new_n949), .A3(new_n950), .A4(new_n425), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n379), .A2(new_n384), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT16), .B1(new_n952), .B2(new_n400), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n369), .B1(new_n408), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n946), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT106), .B(new_n369), .C1(new_n408), .C2(new_n953), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n956), .A2(new_n417), .A3(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n425), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n951), .B1(new_n961), .B2(KEYINPUT37), .ZN(new_n962));
  INV_X1    g0762(.A(new_n959), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n429), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n944), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n961), .A2(KEYINPUT37), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n949), .A2(new_n950), .A3(new_n945), .A4(new_n425), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n944), .B1(new_n429), .B2(new_n963), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n943), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n711), .A2(new_n948), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n964), .A2(KEYINPUT38), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n962), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n425), .B1(new_n367), .B2(new_n398), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n946), .B(KEYINPUT107), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n398), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT37), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n968), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n429), .A2(new_n979), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT38), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n976), .A2(KEYINPUT39), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n972), .A2(KEYINPUT39), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n296), .A2(new_n731), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n973), .B(new_n974), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n778), .A2(new_n464), .A3(new_n793), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n716), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n988), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n465), .A2(new_n770), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n939), .A2(new_n890), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT108), .B1(new_n993), .B2(new_n770), .ZN(new_n994));
  AND4_X1   g0794(.A1(new_n578), .A2(new_n620), .A3(new_n628), .A4(new_n674), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n743), .A2(new_n995), .A3(new_n737), .ZN(new_n996));
  INV_X1    g0796(.A(new_n768), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n766), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT40), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT108), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n999), .A2(new_n890), .A3(new_n939), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(new_n972), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n976), .A2(new_n983), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n999), .A2(new_n890), .A3(new_n939), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT40), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n771), .B1(new_n992), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n992), .B2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n991), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n203), .B2(new_n797), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n991), .A2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n931), .B1(new_n1011), .B2(new_n1012), .ZN(G367));
  OAI221_X1 g0813(.A(new_n871), .B1(new_n207), .B2(new_n455), .C1(new_n873), .C2(new_n233), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n883), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n731), .A2(new_n695), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n682), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n677), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n812), .A2(new_n246), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n855), .A2(new_n309), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(G50), .C2(new_n836), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n273), .B1(new_n910), .B2(new_n839), .C1(new_n825), .C2(new_n248), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n820), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1024), .A2(G58), .B1(G137), .B2(new_n832), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1022), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n852), .A2(G159), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1021), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n850), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n872), .B1(new_n833), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G97), .B2(new_n824), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT46), .B1(new_n1024), .B2(new_n496), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G303), .B2(new_n830), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1030), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n812), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n438), .B1(new_n836), .B2(G283), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n859), .B2(new_n839), .C1(new_n848), .C2(new_n860), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1029), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  OAI221_X1 g0841(.A(new_n1015), .B1(new_n880), .B2(new_n1018), .C1(new_n1041), .C2(new_n807), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n620), .B(new_n628), .C1(new_n624), .C2(new_n737), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n787), .A2(new_n731), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n745), .A2(new_n742), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT45), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n745), .A2(new_n742), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT44), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT44), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1053), .B(new_n1045), .C1(new_n745), .C2(new_n742), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1048), .A2(new_n1049), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n741), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n745), .B1(new_n740), .B2(new_n744), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(new_n736), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n794), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n748), .B(KEYINPUT41), .Z(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n800), .A2(new_n203), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1056), .A2(new_n1045), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT110), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1018), .B(KEYINPUT43), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1045), .A2(new_n743), .A3(new_n744), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT42), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(KEYINPUT109), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT109), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1069), .B2(KEYINPUT42), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n620), .B1(new_n1043), .B2(new_n739), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1069), .A2(KEYINPUT42), .B1(new_n737), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1068), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1077), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1074), .B2(new_n1072), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1078), .A2(KEYINPUT111), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT111), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1080), .B2(new_n1068), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1067), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1067), .A3(new_n1084), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(KEYINPUT112), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT112), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1082), .A2(new_n1088), .A3(new_n1067), .A4(new_n1084), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1065), .A2(new_n1090), .A3(KEYINPUT113), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT113), .B1(new_n1065), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1042), .B1(new_n1091), .B2(new_n1092), .ZN(G387));
  INV_X1    g0893(.A(new_n1059), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1064), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n740), .A2(new_n880), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n750), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n876), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(G107), .B2(new_n207), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n230), .A2(new_n268), .ZN(new_n1100));
  AOI211_X1 g0900(.A(G45), .B(new_n1097), .C1(G68), .C2(G77), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n308), .A2(G50), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n873), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n871), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n883), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n812), .A2(new_n455), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n837), .A2(new_n246), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G50), .C2(new_n830), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n308), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n852), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n833), .A2(new_n309), .B1(new_n248), .B2(new_n820), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n872), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n834), .B2(new_n839), .C1(new_n825), .C2(new_n597), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1116), .B2(new_n1115), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1112), .A2(new_n1114), .A3(new_n1117), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n820), .A2(new_n860), .B1(new_n812), .B2(new_n863), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G317), .A2(new_n830), .B1(new_n901), .B2(G322), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n537), .B2(new_n837), .C1(new_n848), .C2(new_n859), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT48), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT49), .Z(new_n1128));
  OAI221_X1 g0928(.A(new_n872), .B1(new_n825), .B2(new_n552), .C1(new_n833), .C2(new_n857), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1121), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1109), .B1(new_n1130), .B2(new_n806), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1094), .A2(new_n1095), .B1(new_n1096), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1094), .A2(new_n794), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n748), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1094), .A2(new_n794), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(G393));
  OAI221_X1 g0936(.A(new_n871), .B1(new_n597), .B2(new_n207), .C1(new_n873), .C2(new_n243), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n883), .A2(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n855), .A2(new_n859), .B1(new_n1031), .B2(new_n839), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT52), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n833), .A2(new_n856), .B1(new_n863), .B2(new_n820), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n837), .A2(new_n860), .B1(new_n552), .B2(new_n812), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n320), .B1(new_n825), .B2(new_n434), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1140), .B(new_n1144), .C1(new_n537), .C2(new_n848), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n855), .A2(new_n834), .B1(new_n309), .B2(new_n839), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT51), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1037), .A2(G77), .B1(new_n836), .B2(new_n1113), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n838), .C2(new_n848), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n872), .B1(new_n824), .B2(G87), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n246), .B2(new_n820), .C1(new_n910), .C2(new_n833), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT117), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n1145), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1138), .B1(new_n1153), .B2(new_n806), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1045), .B2(new_n880), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1057), .A2(new_n1133), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n748), .B1(new_n1057), .B2(new_n1133), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1155), .B1(new_n1057), .B2(new_n1064), .C1(new_n1156), .C2(new_n1157), .ZN(G390));
  AOI22_X1  g0958(.A1(G132), .A2(new_n830), .B1(new_n901), .B2(G128), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1159), .B1(new_n834), .B2(new_n812), .C1(new_n837), .C2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n820), .A2(new_n309), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n320), .B1(new_n824), .B2(G50), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1165), .C1(new_n1166), .C2(new_n833), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1161), .B(new_n1167), .C1(G137), .C2(new_n852), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n320), .B1(new_n248), .B2(new_n812), .C1(new_n905), .C2(new_n668), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n914), .B1(new_n833), .B2(new_n860), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT121), .Z(new_n1171));
  AOI22_X1  g0971(.A1(G116), .A2(new_n830), .B1(new_n901), .B2(G283), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n597), .B2(new_n837), .C1(new_n848), .C2(new_n439), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n806), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n805), .B1(new_n308), .B2(new_n898), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n986), .B2(new_n868), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n780), .A2(new_n677), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n700), .A2(KEYINPUT26), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n890), .B(new_n737), .C1(new_n688), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n940), .B1(new_n1182), .B2(new_n942), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n987), .B1(new_n976), .B2(new_n983), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT118), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT118), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n987), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n981), .A2(new_n982), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n944), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n971), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n941), .B1(new_n792), .B2(new_n890), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1186), .B(new_n1190), .C1(new_n1191), .C2(new_n940), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1185), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n984), .B(new_n985), .C1(new_n1187), .C2(new_n943), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n999), .A2(G330), .A3(new_n890), .A4(new_n939), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1178), .B1(new_n1198), .B2(new_n1095), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G330), .B(new_n890), .C1(new_n754), .C2(new_n769), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n940), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n893), .A2(new_n942), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n464), .A2(new_n772), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n716), .A3(new_n989), .A4(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(KEYINPUT119), .B(new_n1207), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1195), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n989), .A2(new_n716), .A3(new_n1206), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1201), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1201), .A2(new_n1195), .B1(new_n893), .B2(new_n942), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1208), .A2(new_n748), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1217), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT119), .B1(new_n1220), .B2(new_n1207), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1199), .B1(new_n1219), .B2(new_n1221), .ZN(G378));
  AOI21_X1  g1022(.A(new_n805), .B1(new_n838), .B2(new_n898), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n872), .A2(new_n267), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n824), .A2(G58), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n833), .B2(new_n863), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G77), .C2(new_n1024), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1019), .B1(new_n647), .B2(new_n836), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G107), .A2(new_n830), .B1(new_n901), .B2(G116), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n852), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT58), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT58), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1224), .B(new_n838), .C1(G33), .C2(G41), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n316), .B(new_n267), .C1(new_n825), .C2(new_n834), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n830), .A2(G128), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n820), .B2(new_n1160), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n836), .A2(G137), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n1166), .B2(new_n839), .C1(new_n309), .C2(new_n812), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G132), .C2(new_n852), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT59), .Z(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1236), .B(new_n1243), .C1(G124), .C2(new_n832), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1223), .B1(new_n1246), .B2(new_n807), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n314), .A2(new_n946), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n703), .B2(new_n335), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1249), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n349), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1248), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1252), .A3(new_n1248), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(KEYINPUT123), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1250), .A2(new_n1252), .A3(new_n1248), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1253), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1247), .B1(new_n1260), .B2(new_n868), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n973), .A2(new_n974), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n986), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1187), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1007), .A2(new_n1260), .A3(G330), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n771), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1258), .A2(new_n1253), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1260), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n988), .B(new_n1270), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1261), .B1(new_n1272), .B2(new_n1095), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1212), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1218), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1272), .A3(KEYINPUT57), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n748), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1275), .B2(new_n1272), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(G375));
  NAND2_X1  g1079(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1207), .A2(new_n1062), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n805), .B1(new_n246), .B2(new_n898), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n852), .A2(new_n496), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n863), .A2(new_n855), .B1(new_n837), .B2(new_n439), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1110), .B(new_n1284), .C1(G294), .C2(new_n901), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n850), .A2(G97), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n320), .B1(new_n825), .B2(new_n248), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G303), .B2(new_n832), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n1283), .A2(new_n1285), .A3(new_n1286), .A4(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n850), .A2(G159), .B1(G128), .B2(new_n832), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT124), .Z(new_n1291));
  AOI22_X1  g1091(.A1(G137), .A2(new_n830), .B1(new_n901), .B2(G132), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n309), .B2(new_n837), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n848), .A2(new_n1160), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1225), .B(new_n1118), .C1(new_n838), .C2(new_n812), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1289), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1282), .B1(new_n939), .B2(new_n869), .C1(new_n807), .C2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1215), .B2(new_n1064), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1281), .A2(new_n1300), .ZN(G381));
  INV_X1    g1101(.A(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n919), .ZN(new_n1303));
  OR4_X1    g1103(.A1(G396), .A2(new_n1303), .A3(G393), .A4(G381), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G378), .A2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(KEYINPUT125), .B(new_n1199), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G375), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OR3_X1    g1110(.A1(new_n1304), .A2(new_n1310), .A3(G387), .ZN(G407));
  OAI211_X1 g1111(.A(G407), .B(G213), .C1(G343), .C2(new_n1310), .ZN(G409));
  XOR2_X1   g1112(.A(G393), .B(G396), .Z(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1065), .A2(new_n1090), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT113), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1065), .A2(new_n1090), .A3(KEYINPUT113), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G390), .B1(new_n1319), .B2(new_n1042), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1042), .B(G390), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1302), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(new_n1313), .A3(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n728), .A2(G343), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1275), .A2(new_n1272), .A3(new_n1062), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1273), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1306), .A2(new_n1307), .A3(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G378), .B(new_n1273), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1327), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT60), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1280), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1212), .A2(new_n1215), .A3(KEYINPUT60), .ZN(new_n1335));
  AND4_X1   g1135(.A1(KEYINPUT126), .A2(new_n1334), .A3(new_n748), .A4(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n749), .B1(new_n1333), .B2(new_n1280), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT126), .B1(new_n1337), .B2(new_n1335), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1300), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n919), .ZN(new_n1340));
  OAI211_X1 g1140(.A(G384), .B(new_n1300), .C1(new_n1336), .C2(new_n1338), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1332), .A2(KEYINPUT62), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT62), .B1(new_n1332), .B2(new_n1343), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT127), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1327), .A2(G2897), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1340), .A2(new_n1341), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1327), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1352), .A2(new_n1343), .A3(new_n1353), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT62), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1346), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1326), .B1(new_n1347), .B2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT63), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1326), .B1(new_n1361), .B2(new_n1356), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1332), .A2(KEYINPUT63), .A3(new_n1343), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1362), .A2(new_n1363), .A3(new_n1355), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1360), .A2(new_n1364), .ZN(G405));
  NAND2_X1  g1165(.A1(new_n1308), .A2(G375), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1331), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(new_n1367), .B(new_n1343), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1368), .B(new_n1326), .ZN(G402));
endmodule


