//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT80), .A2(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT80), .A2(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(new_n192), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G107), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT80), .A2(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT80), .A2(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n198), .A2(new_n195), .A3(G107), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n194), .B1(new_n197), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n194), .B(new_n204), .C1(new_n197), .C2(new_n201), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT2), .A2(G113), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT2), .A2(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT2), .A3(G113), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G116), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n212), .B(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n198), .A2(G107), .A3(new_n199), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n200), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n204), .B1(new_n222), .B2(new_n194), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n219), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n193), .B1(G104), .B2(new_n190), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n205), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n214), .A3(G116), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n233), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT84), .B1(new_n231), .B2(new_n234), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n206), .A2(new_n225), .B1(new_n228), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n187), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n240), .B2(KEYINPUT85), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n206), .A2(new_n225), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n228), .A2(new_n239), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n245), .A2(KEYINPUT85), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n242), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n246), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n187), .A3(new_n252), .A4(new_n243), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT64), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT0), .B(G128), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT64), .A2(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT64), .A2(G143), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n256), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT65), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n255), .A2(G143), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(new_n272), .C1(new_n261), .C2(new_n255), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT1), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n272), .B(new_n277), .C1(new_n261), .C2(new_n255), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n262), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G224), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G953), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n248), .A2(new_n253), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n282), .A2(new_n284), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n287), .A2(KEYINPUT7), .B1(new_n240), .B2(new_n241), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n241), .B(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n205), .A2(new_n227), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n235), .A2(new_n230), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n290), .B2(new_n239), .ZN(new_n293));
  INV_X1    g107(.A(new_n284), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n275), .A2(new_n281), .B1(KEYINPUT7), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT86), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n286), .A2(new_n304), .A3(new_n297), .A4(new_n298), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G953), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n307), .A2(G952), .ZN(new_n308));
  INV_X1    g122(.A(G234), .ZN(new_n309));
  INV_X1    g123(.A(G237), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT73), .B(G902), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n307), .B(new_n313), .C1(G234), .C2(G237), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT95), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n321));
  NOR2_X1   g135(.A1(G475), .A2(G902), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n310), .A2(new_n307), .A3(G143), .A4(G214), .ZN(new_n323));
  INV_X1    g137(.A(G214), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n324), .A2(G237), .A3(G953), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT87), .B(new_n323), .C1(new_n261), .C2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(G143), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(KEYINPUT18), .A3(G131), .A4(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(new_n255), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n255), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n323), .A2(KEYINPUT87), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n325), .B2(G143), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n265), .A2(new_n266), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n310), .A2(new_n307), .A3(G214), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT18), .A2(G131), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n329), .B(new_n333), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n326), .A2(G131), .A3(new_n328), .ZN(new_n343));
  AOI21_X1  g157(.A(G131), .B1(new_n326), .B2(new_n328), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G125), .ZN(new_n346));
  OR3_X1    g160(.A1(new_n346), .A2(KEYINPUT16), .A3(G140), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n346), .A2(KEYINPUT16), .A3(G140), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n351));
  OAI211_X1 g165(.A(G146), .B(new_n349), .C1(new_n351), .C2(new_n348), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n330), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(new_n255), .C1(new_n330), .C2(new_n354), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n342), .B1(new_n345), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G113), .B(G122), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(new_n188), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(KEYINPUT89), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n346), .A2(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n348), .B1(new_n366), .B2(new_n347), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n255), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n339), .A2(G131), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n352), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT17), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n360), .B(new_n342), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT89), .B1(new_n358), .B2(new_n361), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n321), .B(new_n322), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT90), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n326), .A2(new_n328), .ZN(new_n380));
  INV_X1    g194(.A(G131), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n370), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n352), .A2(new_n356), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n380), .A2(new_n340), .B1(new_n332), .B2(new_n331), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n329), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n386), .B2(new_n360), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n374), .A3(new_n362), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n321), .A4(new_n322), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n322), .B1(new_n375), .B2(new_n376), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT20), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n378), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT15), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(KEYINPUT15), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G116), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n216), .A2(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(G107), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT91), .B1(new_n258), .B2(G128), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT91), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n276), .A3(G143), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n259), .A2(G128), .A3(new_n260), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT66), .B(G134), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT13), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT13), .B1(new_n336), .B2(G128), .ZN(new_n416));
  OAI21_X1  g230(.A(G134), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT92), .B(G134), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n411), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n190), .B1(new_n402), .B2(KEYINPUT14), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(new_n404), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(G953), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT93), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n413), .ZN(new_n432));
  INV_X1    g246(.A(new_n420), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n410), .A2(new_n414), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n336), .A2(KEYINPUT13), .A3(G128), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n409), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT92), .B1(new_n436), .B2(G134), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n423), .A2(new_n425), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT93), .A4(new_n430), .ZN(new_n440));
  INV_X1    g254(.A(new_n430), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n421), .B2(new_n426), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n313), .B(new_n400), .C1(new_n431), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n439), .A3(new_n430), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n442), .A3(new_n440), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n400), .B1(new_n449), .B2(new_n313), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n342), .B1(new_n372), .B2(new_n373), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n361), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n374), .ZN(new_n454));
  INV_X1    g268(.A(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G475), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n393), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n272), .B1(new_n261), .B2(new_n255), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT1), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n261), .B2(new_n255), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n464), .B2(new_n276), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n336), .A2(G146), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(KEYINPUT82), .A3(new_n272), .A4(new_n277), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n278), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n461), .B1(new_n471), .B2(new_n290), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n273), .B1(new_n269), .B2(KEYINPUT65), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n254), .B(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n202), .A2(new_n224), .A3(G101), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n205), .A2(KEYINPUT4), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n223), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n205), .A2(KEYINPUT10), .A3(new_n280), .A4(new_n227), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT11), .ZN(new_n481));
  INV_X1    g295(.A(G134), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G134), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n485), .A3(G137), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n482), .A2(G137), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n481), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n485), .ZN(new_n490));
  INV_X1    g304(.A(G137), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT11), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n481), .B1(new_n411), .B2(G137), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n411), .B2(G137), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n381), .B(new_n494), .C1(new_n495), .C2(new_n481), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n480), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n493), .A2(new_n496), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n472), .A2(new_n478), .A3(new_n499), .A4(new_n479), .ZN(new_n500));
  XNOR2_X1  g314(.A(G110), .B(G140), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n307), .A2(G227), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n280), .B1(new_n205), .B2(new_n227), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n228), .B2(new_n470), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n497), .A2(KEYINPUT83), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT12), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n510));
  INV_X1    g324(.A(new_n508), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n471), .A2(new_n290), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n511), .C1(new_n512), .C2(new_n506), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n500), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n498), .A2(new_n505), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  OAI21_X1  g329(.A(G469), .B1(new_n515), .B2(G902), .ZN(new_n516));
  INV_X1    g330(.A(G469), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n504), .A2(new_n509), .A3(new_n500), .A4(new_n513), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n504), .B1(new_n498), .B2(new_n500), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n517), .B(new_n313), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n460), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  AND4_X1   g335(.A1(new_n306), .A2(new_n320), .A3(new_n458), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n310), .A2(new_n307), .A3(G210), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n524), .B(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n527), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(G101), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n538));
  AOI21_X1  g352(.A(G137), .B1(new_n483), .B2(new_n485), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n491), .A2(G134), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n538), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n540), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n411), .B2(G137), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n538), .B1(new_n544), .B2(G131), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n496), .B(new_n280), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n499), .B2(new_n274), .ZN(new_n547));
  INV_X1    g361(.A(new_n219), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n475), .A2(new_n497), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n219), .A3(new_n546), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n537), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n542), .A2(new_n545), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n496), .A2(new_n280), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(new_n554), .B1(new_n475), .B2(new_n497), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT28), .B1(new_n555), .B2(new_n219), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n536), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n550), .A2(new_n558), .A3(new_n546), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n550), .B2(new_n546), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n548), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n551), .A2(new_n535), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n547), .A2(KEYINPUT30), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n550), .A2(new_n558), .A3(new_n546), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n219), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT31), .B1(new_n569), .B2(new_n563), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n561), .A2(new_n564), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT32), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n569), .A2(KEYINPUT31), .A3(new_n563), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n550), .A2(new_n219), .A3(new_n546), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n219), .B1(new_n550), .B2(new_n546), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT28), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n551), .A2(new_n537), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n535), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT72), .B1(new_n573), .B2(KEYINPUT31), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n571), .B(new_n562), .C1(new_n561), .C2(new_n564), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n576), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n582), .A2(KEYINPUT29), .A3(new_n535), .A4(new_n583), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n313), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n536), .B1(new_n569), .B2(new_n580), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n549), .A2(new_n551), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n556), .B1(new_n595), .B2(KEYINPUT28), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT29), .B1(new_n596), .B2(new_n535), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n593), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G472), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n592), .A2(new_n313), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT29), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n582), .A2(new_n535), .A3(new_n583), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n594), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n599), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT74), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n578), .A2(new_n590), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n429), .B1(new_n313), .B2(G234), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n214), .A2(G128), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT23), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT76), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n214), .A2(G128), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(KEYINPUT23), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n615), .B2(new_n610), .ZN(new_n616));
  INV_X1    g430(.A(G110), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n276), .B2(G119), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n214), .A2(KEYINPUT75), .A3(G128), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n276), .A2(G119), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT24), .B(G110), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n616), .A2(new_n617), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n352), .B2(new_n369), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n332), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n367), .A2(new_n368), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(G146), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT23), .B1(new_n276), .B2(G119), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n610), .B1(new_n632), .B2(KEYINPUT76), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n622), .A2(new_n613), .A3(KEYINPUT23), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n617), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT78), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(KEYINPUT78), .A3(new_n352), .A4(new_n332), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n627), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT22), .B(G137), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n636), .A2(new_n352), .A3(new_n332), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT78), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n626), .B1(new_n647), .B2(new_n638), .ZN(new_n648));
  INV_X1    g462(.A(new_n643), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n313), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT25), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n644), .A2(new_n650), .A3(KEYINPUT25), .A4(new_n313), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n609), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n648), .A2(new_n649), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n643), .B(new_n626), .C1(new_n647), .C2(new_n638), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n608), .A2(G902), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT79), .B1(new_n607), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n577), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n589), .B1(new_n588), .B2(new_n576), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n605), .A2(KEYINPUT74), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n591), .B(new_n599), .C1(new_n601), .C2(new_n604), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n666), .A2(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT79), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n663), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n523), .B1(new_n665), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n204), .ZN(G3));
  NAND2_X1  g488(.A1(new_n505), .A2(new_n498), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n514), .A2(new_n503), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(G469), .ZN(new_n677));
  NAND2_X1  g491(.A1(G469), .A2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n520), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n663), .A3(new_n459), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n599), .B1(new_n588), .B2(new_n313), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n575), .A2(new_n577), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n317), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n286), .A2(new_n297), .A3(new_n298), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n298), .B1(new_n286), .B2(new_n297), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n684), .B(new_n318), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n393), .A2(new_n457), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n442), .A2(new_n446), .A3(KEYINPUT33), .ZN(new_n689));
  INV_X1    g503(.A(new_n313), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n394), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n431), .A2(new_n443), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n689), .B(new_n691), .C1(new_n692), .C2(KEYINPUT33), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n313), .B1(new_n431), .B2(new_n443), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n394), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT34), .B(G104), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G6));
  INV_X1    g516(.A(new_n377), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n321), .B1(new_n388), .B2(new_n322), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n457), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n451), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n684), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n318), .B1(new_n685), .B2(new_n686), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n683), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT35), .B(G107), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G9));
  INV_X1    g526(.A(KEYINPUT98), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n575), .B2(new_n690), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n588), .A2(new_n576), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT25), .B1(new_n658), .B2(new_n313), .ZN(new_n717));
  INV_X1    g531(.A(new_n654), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n608), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT97), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n643), .A2(KEYINPUT36), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n648), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n648), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n660), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n725), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT97), .B1(new_n655), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n713), .B1(new_n716), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n720), .B1(new_n719), .B2(new_n725), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n655), .A2(new_n727), .A3(KEYINPUT97), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT98), .A3(new_n715), .A4(new_n714), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n522), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT37), .B(G110), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G12));
  NAND3_X1  g551(.A1(new_n670), .A2(new_n521), .A3(new_n733), .ZN(new_n738));
  INV_X1    g552(.A(G900), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n314), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n311), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT99), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n706), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT100), .B1(new_n743), .B2(new_n708), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n319), .B1(new_n303), .B2(new_n299), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT100), .ZN(new_n746));
  INV_X1    g560(.A(new_n742), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n705), .A2(new_n451), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n276), .ZN(G30));
  XNOR2_X1  g566(.A(new_n742), .B(KEYINPUT39), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n521), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT40), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n306), .B(KEYINPUT38), .Z(new_n756));
  AOI21_X1  g570(.A(new_n536), .B1(new_n561), .B2(new_n551), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n455), .B1(new_n595), .B2(new_n535), .ZN(new_n758));
  OAI21_X1  g572(.A(G472), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n666), .B2(new_n667), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n655), .A2(new_n727), .ZN(new_n761));
  INV_X1    g575(.A(new_n688), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n451), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n318), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n755), .A2(new_n756), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n261), .ZN(G45));
  NAND3_X1  g580(.A1(new_n688), .A2(new_n696), .A3(new_n742), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n708), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n670), .A2(new_n521), .A3(new_n733), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G146), .ZN(G48));
  OAI21_X1  g584(.A(new_n313), .B1(new_n518), .B2(new_n519), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(G469), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n459), .A3(new_n520), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n670), .A2(new_n663), .A3(new_n698), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n578), .A2(new_n590), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n600), .A2(new_n606), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n664), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT101), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n780), .A3(new_n698), .A4(new_n774), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT41), .B(G113), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G15));
  NAND4_X1  g598(.A1(new_n670), .A2(new_n709), .A3(new_n663), .A4(new_n774), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT102), .B(G116), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G18));
  NAND4_X1  g601(.A1(new_n393), .A2(new_n451), .A3(new_n684), .A4(new_n457), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n708), .A2(new_n773), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n670), .A2(new_n789), .A3(new_n733), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G119), .ZN(G21));
  NAND3_X1  g605(.A1(new_n557), .A2(new_n570), .A3(new_n565), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n576), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT103), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT103), .A3(new_n576), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n681), .A3(new_n664), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n694), .A2(new_n399), .ZN(new_n799));
  AOI221_X4 g613(.A(KEYINPUT104), .B1(new_n799), .B2(new_n444), .C1(new_n393), .C2(new_n457), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT104), .ZN(new_n801));
  INV_X1    g615(.A(new_n451), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n688), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n708), .A2(new_n773), .A3(new_n317), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n798), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT105), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT105), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n798), .A2(new_n804), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G122), .ZN(G24));
  NOR3_X1   g625(.A1(new_n797), .A2(new_n681), .A3(new_n761), .ZN(new_n812));
  AOI221_X4 g626(.A(new_n747), .B1(new_n693), .B2(new_n695), .C1(new_n393), .C2(new_n457), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n708), .A2(new_n773), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G125), .ZN(G27));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n666), .B2(new_n667), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n578), .A2(KEYINPUT108), .A3(new_n590), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n778), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n300), .A2(new_n303), .A3(new_n305), .A4(new_n318), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n678), .B(KEYINPUT106), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n520), .A2(new_n677), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n459), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT42), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n821), .A2(new_n767), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n826), .A3(new_n663), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n820), .A2(new_n826), .A3(new_n829), .A4(new_n663), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n821), .A2(new_n824), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n779), .A2(new_n813), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n828), .A2(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n381), .ZN(G33));
  NAND3_X1  g649(.A1(new_n779), .A2(new_n748), .A3(new_n831), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G134), .ZN(G36));
  AOI21_X1  g651(.A(new_n688), .B1(new_n695), .B2(new_n693), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT43), .ZN(new_n839));
  INV_X1    g653(.A(new_n761), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n839), .A2(new_n716), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n821), .B1(new_n841), .B2(KEYINPUT44), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(KEYINPUT44), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g657(.A(G469), .B1(new_n515), .B2(KEYINPUT45), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(KEYINPUT45), .B2(new_n515), .ZN(new_n845));
  INV_X1    g659(.A(new_n822), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT46), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n847), .B2(KEYINPUT46), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(KEYINPUT46), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n520), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n459), .ZN(new_n853));
  INV_X1    g667(.A(new_n753), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n853), .A2(KEYINPUT111), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT111), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n843), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(new_n491), .ZN(G39));
  INV_X1    g672(.A(KEYINPUT47), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(KEYINPUT47), .A3(new_n459), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n670), .A2(new_n663), .A3(new_n767), .A4(new_n821), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n363), .ZN(G42));
  AND2_X1   g679(.A1(new_n839), .A2(new_n312), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n798), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n814), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT120), .Z(new_n869));
  AOI22_X1  g683(.A1(new_n777), .A2(new_n817), .B1(new_n600), .B2(new_n606), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n664), .B1(new_n870), .B2(new_n819), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n821), .A2(new_n773), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT48), .ZN(new_n874));
  INV_X1    g688(.A(new_n760), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n663), .A3(new_n312), .A4(new_n872), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(new_n697), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n869), .A2(new_n308), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n867), .A2(new_n319), .A3(new_n756), .A4(new_n774), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT50), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n821), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n772), .A2(new_n520), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n459), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n882), .B(new_n867), .C1(new_n862), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n866), .A2(new_n812), .A3(new_n872), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n876), .A2(new_n688), .A3(new_n696), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n881), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n889), .B2(new_n888), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(new_n796), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT103), .B1(new_n792), .B2(new_n576), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n714), .A3(new_n840), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n774), .A2(new_n745), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n767), .ZN(new_n898));
  INV_X1    g712(.A(new_n521), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n607), .A2(new_n899), .A3(new_n729), .ZN(new_n900));
  INV_X1    g714(.A(new_n750), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n459), .A2(new_n823), .A3(new_n761), .A4(new_n742), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n804), .A2(new_n760), .A3(new_n903), .A4(new_n745), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n769), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n815), .B1(new_n738), .B2(new_n750), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT118), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT118), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n769), .A3(new_n904), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n912), .B2(KEYINPUT52), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n832), .A2(new_n833), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n829), .B1(new_n871), .B2(new_n826), .ZN(new_n915));
  INV_X1    g729(.A(new_n830), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n812), .A2(new_n813), .A3(new_n831), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n836), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n729), .B1(new_n777), .B2(new_n778), .ZN(new_n920));
  AOI22_X1  g734(.A1(new_n392), .A2(new_n377), .B1(G475), .B2(new_n456), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n451), .A3(new_n922), .A4(new_n742), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n799), .A2(new_n444), .A3(new_n742), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT114), .B1(new_n705), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n882), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT115), .B1(new_n929), .B2(new_n821), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n920), .A2(new_n928), .A3(new_n521), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n900), .A2(KEYINPUT116), .A3(new_n930), .A4(new_n928), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n919), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n917), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n306), .A2(new_n320), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n688), .A2(new_n451), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n683), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n735), .A2(new_n785), .A3(new_n790), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n673), .ZN(new_n941));
  AOI22_X1  g755(.A1(new_n781), .A2(new_n776), .B1(new_n807), .B2(new_n809), .ZN(new_n942));
  INV_X1    g756(.A(new_n697), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT113), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT113), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n683), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n942), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n936), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n913), .A2(new_n950), .A3(KEYINPUT53), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT119), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n769), .A2(new_n904), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT52), .B1(new_n909), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n907), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n907), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT117), .B1(new_n936), .B2(new_n949), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n782), .A2(new_n810), .A3(new_n948), .ZN(new_n959));
  AOI211_X1 g773(.A(KEYINPUT79), .B(new_n664), .C1(new_n777), .C2(new_n778), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n671), .B1(new_n670), .B2(new_n663), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n522), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n938), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n716), .A2(new_n963), .A3(new_n680), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n964), .A2(new_n937), .B1(new_n920), .B2(new_n789), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n962), .A2(new_n735), .A3(new_n785), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT117), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n917), .A4(new_n935), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n957), .B1(new_n958), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n892), .B(new_n951), .C1(new_n970), .C2(KEYINPUT53), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n958), .A2(new_n969), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT53), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n913), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n973), .B2(new_n970), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n975), .B2(new_n892), .ZN(new_n976));
  OAI22_X1  g790(.A1(new_n891), .A2(new_n976), .B1(G952), .B2(G953), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n883), .A2(KEYINPUT49), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n883), .A2(KEYINPUT49), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n663), .A2(new_n318), .A3(new_n459), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n756), .A2(new_n875), .A3(new_n838), .A4(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n977), .A2(new_n983), .ZN(G75));
  INV_X1    g798(.A(KEYINPUT56), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n248), .A2(new_n253), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n285), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT55), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n955), .A2(new_n956), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT53), .B1(new_n972), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n951), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n313), .A2(new_n298), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n985), .B(new_n989), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n307), .A2(KEYINPUT122), .A3(G952), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT122), .B1(new_n307), .B2(G952), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT121), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n933), .A2(new_n934), .ZN(new_n1003));
  INV_X1    g817(.A(new_n919), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1005), .A2(new_n834), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n968), .B1(new_n1006), .B2(new_n967), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n936), .A2(new_n949), .A3(KEYINPUT117), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n990), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n973), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n951), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT56), .B1(new_n1011), .B2(new_n994), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1002), .B1(new_n1012), .B2(new_n989), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n985), .B1(new_n993), .B2(new_n995), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(KEYINPUT121), .A3(new_n988), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1001), .B1(new_n1013), .B2(new_n1015), .ZN(G51));
  XOR2_X1   g830(.A(new_n822), .B(KEYINPUT57), .Z(new_n1017));
  AOI21_X1  g831(.A(new_n892), .B1(new_n1010), .B2(new_n951), .ZN(new_n1018));
  INV_X1    g832(.A(new_n971), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n518), .A2(new_n519), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1011), .A2(new_n690), .A3(new_n845), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n999), .B1(new_n1022), .B2(new_n1023), .ZN(G54));
  INV_X1    g838(.A(KEYINPUT124), .ZN(new_n1025));
  AND2_X1   g839(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n690), .B(new_n1026), .C1(new_n991), .C2(new_n992), .ZN(new_n1027));
  INV_X1    g841(.A(new_n388), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n388), .A2(new_n1026), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n690), .B(new_n1030), .C1(new_n991), .C2(new_n992), .ZN(new_n1031));
  INV_X1    g845(.A(new_n999), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1025), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1035), .A2(KEYINPUT124), .A3(new_n1032), .A4(new_n1031), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(G60));
  OAI21_X1  g851(.A(new_n689), .B1(new_n692), .B2(KEYINPUT33), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G478), .A2(G902), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT59), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1039), .B1(new_n976), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1000), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1044));
  OAI21_X1  g858(.A(KEYINPUT54), .B1(new_n991), .B2(new_n992), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n1045), .B2(new_n971), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(G63));
  NAND2_X1  g861(.A1(G217), .A2(G902), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT125), .Z(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT60), .Z(new_n1050));
  OAI211_X1 g864(.A(new_n724), .B(new_n1050), .C1(new_n991), .C2(new_n992), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1050), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n1010), .B2(new_n951), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n1000), .B(new_n1051), .C1(new_n1053), .C2(new_n658), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT61), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n659), .B1(new_n993), .B2(new_n1052), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1057), .A2(KEYINPUT61), .A3(new_n1000), .A4(new_n1051), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1056), .A2(new_n1058), .ZN(G66));
  XNOR2_X1  g873(.A(new_n949), .B(KEYINPUT126), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(new_n307), .ZN(new_n1061));
  OAI21_X1  g875(.A(G953), .B1(new_n316), .B2(new_n283), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n986), .B1(G898), .B2(new_n307), .ZN(new_n1064));
  XNOR2_X1  g878(.A(new_n1064), .B(KEYINPUT127), .ZN(new_n1065));
  XNOR2_X1  g879(.A(new_n1063), .B(new_n1065), .ZN(G69));
  NOR2_X1   g880(.A1(new_n857), .A2(new_n864), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n910), .A2(new_n765), .A3(new_n769), .A4(new_n911), .ZN(new_n1068));
  OR2_X1    g882(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1070));
  AOI211_X1 g884(.A(new_n821), .B(new_n754), .C1(new_n697), .C2(new_n963), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1071), .B1(new_n960), .B2(new_n961), .ZN(new_n1072));
  NAND4_X1  g886(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1073), .A2(new_n307), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n559), .A2(new_n560), .ZN(new_n1075));
  OAI21_X1  g889(.A(new_n355), .B1(new_n330), .B2(new_n354), .ZN(new_n1076));
  XOR2_X1   g890(.A(new_n1075), .B(new_n1076), .Z(new_n1077));
  NAND2_X1  g891(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g892(.A(new_n1077), .B1(G900), .B2(G953), .ZN(new_n1079));
  NAND3_X1  g893(.A1(new_n871), .A2(new_n745), .A3(new_n804), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n1080), .B1(new_n855), .B2(new_n856), .ZN(new_n1081));
  NAND3_X1  g895(.A1(new_n910), .A2(new_n769), .A3(new_n911), .ZN(new_n1082));
  NOR2_X1   g896(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g897(.A1(new_n1067), .A2(new_n1083), .A3(new_n917), .A4(new_n836), .ZN(new_n1084));
  OAI21_X1  g898(.A(new_n1079), .B1(new_n1084), .B2(G953), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g900(.A(new_n307), .B1(G227), .B2(G900), .ZN(new_n1087));
  NAND2_X1  g901(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g902(.A(new_n1087), .ZN(new_n1089));
  NAND3_X1  g903(.A1(new_n1078), .A2(new_n1089), .A3(new_n1085), .ZN(new_n1090));
  NAND2_X1  g904(.A1(new_n1088), .A2(new_n1090), .ZN(G72));
  NAND2_X1  g905(.A1(G472), .A2(G902), .ZN(new_n1092));
  XOR2_X1   g906(.A(new_n1092), .B(KEYINPUT63), .Z(new_n1093));
  OAI21_X1  g907(.A(new_n1093), .B1(new_n1084), .B2(new_n1060), .ZN(new_n1094));
  NOR3_X1   g908(.A1(new_n569), .A2(new_n535), .A3(new_n580), .ZN(new_n1095));
  AOI21_X1  g909(.A(new_n999), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g910(.A(new_n757), .ZN(new_n1097));
  NAND2_X1  g911(.A1(new_n1097), .A2(new_n1093), .ZN(new_n1098));
  OR3_X1    g912(.A1(new_n975), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g913(.A(new_n1093), .B1(new_n1073), .B2(new_n1060), .ZN(new_n1100));
  NAND2_X1  g914(.A1(new_n1100), .A2(new_n757), .ZN(new_n1101));
  AND3_X1   g915(.A1(new_n1096), .A2(new_n1099), .A3(new_n1101), .ZN(G57));
endmodule


