//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n217), .A2(new_n218), .B1(new_n206), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n216), .B(new_n220), .C1(G116), .C2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G50), .A2(G226), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n207), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(KEYINPUT65), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n235), .A2(G1), .A3(G13), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G20), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g0040(.A(G50), .B1(G58), .B2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  AOI211_X1 g0042(.A(new_n213), .B(new_n232), .C1(new_n240), .C2(new_n242), .ZN(G361));
  XOR2_X1   g0043(.A(G226), .B(G232), .Z(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G250), .B(G257), .Z(new_n249));
  XNOR2_X1  g0049(.A(G264), .B(G270), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G358));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT67), .B(G107), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(G68), .B(G77), .Z(new_n257));
  XOR2_X1   g0057(.A(G50), .B(G58), .Z(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n263), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(new_n234), .A4(new_n236), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(G20), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n265), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n239), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(G20), .B2(new_n203), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n272), .B1(G50), .B2(new_n273), .C1(new_n274), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT9), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G41), .A2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n270), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT68), .B(G1), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(G226), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n286), .A2(G1), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n237), .A2(new_n291), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT3), .B(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G222), .A2(G1698), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G223), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n301), .B(new_n306), .C1(G77), .C2(new_n302), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n296), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n282), .A2(new_n283), .ZN(new_n310));
  INV_X1    g0110(.A(new_n308), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G190), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n284), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n282), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n290), .A2(G238), .A3(new_n295), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n225), .A2(G1698), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G226), .B2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n298), .B1(new_n301), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n322), .A2(new_n323), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n323), .B1(new_n322), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n334), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(G169), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(G179), .A3(new_n334), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n228), .A2(G20), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n345), .B1(new_n276), .B2(new_n217), .C1(new_n279), .C2(new_n202), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n265), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT72), .B(KEYINPUT11), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n271), .A2(G68), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT12), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n273), .B2(G68), .ZN(new_n352));
  INV_X1    g0152(.A(new_n273), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(KEYINPUT12), .A3(new_n228), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n340), .B2(G200), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n339), .A2(G190), .A3(new_n334), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n344), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n271), .A2(G77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G20), .A2(G77), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n362), .B1(new_n275), .B2(new_n279), .C1(new_n276), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n265), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n353), .A2(new_n217), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n302), .A2(G232), .A3(new_n304), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n302), .A2(G238), .A3(G1698), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(new_n207), .C2(new_n302), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n298), .B1(new_n371), .B2(new_n301), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n290), .A2(G244), .A3(new_n295), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  OAI211_X1 g0175(.A(KEYINPUT71), .B(new_n368), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(G190), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n372), .B2(new_n373), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n367), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n321), .A2(new_n360), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT73), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n330), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n329), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n386));
  OR2_X1    g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n304), .A2(G226), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n301), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n299), .B1(new_n294), .B2(new_n225), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n300), .B1(new_n389), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n375), .B1(new_n397), .B2(new_n393), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(KEYINPUT75), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n392), .A2(new_n394), .A3(new_n400), .A4(new_n395), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT76), .B1(new_n399), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n224), .A2(new_n228), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n201), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n278), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(KEYINPUT7), .B(G20), .C1(new_n385), .C2(new_n386), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT16), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n302), .B2(G20), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n239), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n228), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n408), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n265), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT74), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n273), .A2(new_n275), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n271), .B2(new_n275), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT74), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n414), .A2(new_n425), .A3(new_n265), .A4(new_n420), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n383), .B1(new_n404), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n399), .A2(new_n401), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n401), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n392), .A2(new_n394), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G169), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n315), .B2(new_n437), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT18), .B1(new_n427), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n374), .A2(new_n315), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n372), .A2(new_n373), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n317), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n367), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n382), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n219), .A2(new_n304), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n226), .A2(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n385), .A2(new_n386), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n331), .A2(G303), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n300), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n267), .B2(new_n269), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n458), .A2(G270), .A3(new_n292), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n456), .A2(G274), .A3(new_n292), .A4(new_n457), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR4_X1   g0261(.A1(new_n454), .A2(new_n459), .A3(new_n315), .A4(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n454), .A2(new_n459), .A3(new_n461), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n317), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(KEYINPUT21), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n239), .C1(G33), .C2(new_n206), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT79), .B(G116), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n265), .B(new_n467), .C1(new_n239), .C2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n270), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n274), .A2(new_n273), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(new_n273), .B2(new_n468), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT82), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n454), .A2(new_n461), .ZN(new_n477));
  INV_X1    g0277(.A(new_n459), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT21), .A3(G169), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n463), .A2(G179), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  INV_X1    g0283(.A(new_n475), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n479), .B(G169), .C1(new_n470), .C2(new_n474), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n463), .A2(G190), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n475), .B(new_n489), .C1(new_n375), .C2(new_n463), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n476), .A2(new_n485), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n472), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G87), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n385), .A2(new_n239), .A3(G68), .A4(new_n386), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n239), .B1(new_n324), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G87), .B2(new_n208), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n276), .B2(new_n206), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(new_n265), .B1(new_n353), .B2(new_n363), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n229), .A2(new_n304), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n218), .A2(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n385), .A2(new_n386), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n468), .A2(G33), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n300), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n270), .A2(G45), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n285), .B1(new_n508), .B2(new_n215), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n270), .A2(G45), .A3(new_n297), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n502), .B(new_n512), .C1(new_n375), .C2(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n500), .A2(new_n265), .ZN(new_n515));
  INV_X1    g0315(.A(new_n363), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n274), .A2(new_n273), .A3(new_n516), .A4(new_n471), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n353), .A2(new_n363), .ZN(new_n518));
  AND4_X1   g0318(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n514), .B1(new_n501), .B2(new_n517), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n519), .A2(new_n520), .B1(G169), .B2(new_n511), .ZN(new_n521));
  INV_X1    g0321(.A(new_n507), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n315), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT80), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n513), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n219), .B(new_n285), .C1(new_n456), .C2(new_n457), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT78), .B1(new_n527), .B2(new_n461), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n458), .A2(G257), .A3(new_n292), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(new_n460), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n385), .A2(G244), .A3(new_n304), .A4(new_n386), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n328), .A2(new_n330), .A3(G250), .A4(G1698), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT4), .A2(G244), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n328), .A2(new_n330), .A3(new_n537), .A4(new_n304), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n538), .A3(new_n466), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n300), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n317), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n472), .A2(new_n206), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n273), .A2(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n417), .A2(new_n418), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n279), .A2(new_n217), .ZN(new_n548));
  OR2_X1    g0348(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT6), .A2(G107), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(new_n208), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n553));
  INV_X1    g0353(.A(new_n550), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(G20), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n543), .B(new_n545), .C1(new_n559), .C2(new_n274), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n535), .A2(new_n539), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n301), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(new_n315), .A3(new_n528), .A4(new_n531), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n541), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n274), .B1(new_n547), .B2(new_n558), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n542), .A3(new_n544), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(G190), .A3(new_n528), .A4(new_n531), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n529), .A2(new_n530), .A3(new_n460), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n530), .B1(new_n529), .B2(new_n460), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n568), .A2(new_n540), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n566), .B(new_n567), .C1(new_n570), .C2(new_n375), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n526), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n385), .A2(KEYINPUT22), .A3(G87), .A4(new_n386), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n506), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n239), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n331), .A2(G20), .A3(new_n214), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n239), .A2(G107), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n579), .B(KEYINPUT23), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n576), .A2(KEYINPUT24), .A3(new_n578), .A4(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n265), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n493), .A2(G107), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n273), .A2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n215), .A2(new_n304), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n219), .A2(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n385), .A2(new_n386), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n301), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n458), .A2(G264), .A3(new_n292), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT83), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n300), .B1(new_n592), .B2(new_n593), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n226), .B(new_n285), .C1(new_n456), .C2(new_n457), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT83), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n460), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n598), .A2(new_n599), .A3(new_n461), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n602), .A2(new_n315), .B1(new_n317), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(KEYINPUT84), .A3(new_n375), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT84), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n596), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n600), .B1(new_n598), .B2(new_n599), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n461), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n612), .B2(G200), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n603), .A2(new_n395), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n606), .B1(new_n607), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n449), .A2(new_n492), .A3(new_n573), .A4(new_n616), .ZN(G372));
  AOI22_X1  g0417(.A1(new_n482), .A2(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n572), .B1(new_n605), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT85), .B1(new_n509), .B2(new_n510), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n215), .B1(new_n293), .B2(new_n455), .ZN(new_n621));
  AND4_X1   g0421(.A1(KEYINPUT85), .A2(new_n621), .A3(new_n292), .A4(new_n510), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n522), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n317), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n524), .B(new_n624), .C1(new_n519), .C2(new_n520), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(G200), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n502), .A3(new_n512), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n615), .B2(new_n607), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT86), .B1(new_n619), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n625), .ZN(new_n632));
  XNOR2_X1  g0432(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OR3_X1    g0434(.A1(new_n526), .A2(new_n564), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n564), .A2(KEYINPUT87), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n541), .A2(new_n560), .A3(new_n638), .A4(new_n563), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n640), .B2(new_n628), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n632), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n619), .A2(new_n629), .A3(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n631), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n449), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n319), .ZN(new_n646));
  INV_X1    g0446(.A(new_n442), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n358), .A2(new_n359), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n344), .A2(new_n357), .ZN(new_n649));
  INV_X1    g0449(.A(new_n447), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n651), .B2(new_n436), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n652), .B2(new_n314), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G20), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n293), .A2(new_n657), .A3(KEYINPUT27), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT27), .B1(new_n293), .B2(new_n657), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(G213), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n484), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  INV_X1    g0464(.A(new_n618), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT90), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(KEYINPUT90), .A3(new_n665), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n668), .B(new_n669), .C1(new_n491), .C2(new_n664), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n662), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n616), .B1(new_n607), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n606), .A2(new_n662), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n476), .A2(new_n485), .A3(new_n488), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n616), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n662), .B(KEYINPUT91), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n606), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n675), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n211), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n685), .A2(new_n687), .A3(new_n266), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n690));
  INV_X1    g0490(.A(new_n685), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n689), .B(new_n690), .C1(new_n241), .C2(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n616), .A2(new_n492), .A3(new_n573), .A4(new_n680), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n570), .A2(new_n462), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n511), .B1(new_n597), .B2(new_n601), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n568), .A2(new_n569), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n463), .B1(new_n700), .B2(new_n562), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n315), .A3(new_n602), .A4(new_n623), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n522), .A2(new_n523), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n610), .B2(new_n611), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n570), .A3(KEYINPUT30), .A4(new_n462), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n695), .B1(new_n707), .B2(new_n672), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n699), .A2(new_n702), .A3(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT93), .B1(new_n699), .B2(new_n702), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT31), .B(new_n679), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n694), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n625), .A2(new_n627), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT26), .A3(new_n637), .A4(new_n639), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n634), .B1(new_n526), .B2(new_n564), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n632), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n572), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n629), .B(new_n719), .C1(new_n676), .C2(new_n606), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT94), .B1(new_n721), .B2(new_n672), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT94), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n723), .B(new_n662), .C1(new_n718), .C2(new_n720), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT29), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n644), .A2(new_n680), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n714), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n693), .B1(new_n729), .B2(G1), .ZN(G364));
  OR2_X1    g0530(.A1(new_n670), .A2(G330), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n266), .B1(new_n656), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n685), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n671), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(G20), .A2(G179), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n737), .A2(new_n395), .A3(G200), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  INV_X1    g0539(.A(new_n737), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n739), .A2(G58), .B1(G77), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT97), .Z(new_n745));
  NOR3_X1   g0545(.A1(new_n395), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n239), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n239), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(G97), .B1(new_n751), .B2(G87), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n395), .A3(G200), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n207), .B2(new_n753), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n737), .A2(new_n375), .A3(KEYINPUT98), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT98), .B1(new_n737), .B2(new_n375), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n395), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n331), .B(new_n754), .C1(G50), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n395), .A3(new_n756), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n749), .A2(new_n741), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G159), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n761), .A2(G68), .B1(KEYINPUT32), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n745), .A2(new_n759), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n764), .A2(KEYINPUT32), .ZN(new_n767));
  INV_X1    g0567(.A(new_n758), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n747), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  INV_X1    g0574(.A(new_n753), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n761), .A2(new_n774), .B1(G283), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n331), .B1(new_n750), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n738), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n779), .A2(new_n780), .B1(new_n742), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n778), .B(new_n782), .C1(G329), .C2(new_n763), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n773), .A2(new_n776), .A3(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n766), .A2(new_n767), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n237), .B1(new_n239), .B2(G169), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n385), .A2(new_n386), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n684), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n259), .B2(G45), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n241), .ZN(new_n798));
  NAND3_X1  g0598(.A1(G355), .A2(new_n302), .A3(new_n211), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G116), .C2(new_n211), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n785), .A2(new_n788), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n791), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n734), .B(new_n801), .C1(new_n670), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n736), .A2(new_n803), .ZN(G396));
  AND3_X1   g0604(.A1(new_n619), .A2(new_n629), .A3(KEYINPUT86), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n630), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n679), .B1(new_n806), .B2(new_n642), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT101), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n447), .A2(new_n662), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n367), .A2(new_n662), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n381), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n810), .C1(new_n812), .C2(new_n650), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n650), .B1(new_n381), .B2(new_n811), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT101), .B1(new_n814), .B2(new_n809), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT102), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n813), .A2(new_n815), .A3(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n807), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n714), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n735), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n468), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n770), .A2(new_n779), .B1(new_n828), .B2(new_n742), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n760), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G303), .C2(new_n758), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n751), .A2(G107), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n753), .A2(new_n214), .B1(new_n762), .B2(new_n781), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n302), .B1(new_n834), .B2(KEYINPUT100), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT100), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G97), .B2(new_n748), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G137), .A2(new_n758), .B1(new_n761), .B2(G150), .ZN(new_n839));
  INV_X1    g0639(.A(G159), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n742), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G143), .B2(new_n739), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G132), .B2(new_n763), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n775), .A2(G68), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n748), .A2(G58), .B1(new_n751), .B2(G50), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n838), .B1(new_n847), .B2(new_n793), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n788), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n816), .A2(new_n789), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n788), .A2(new_n789), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n217), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n734), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n827), .A2(new_n853), .ZN(G384));
  INV_X1    g0654(.A(new_n649), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n662), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n416), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n265), .A3(new_n414), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n859), .A2(new_n424), .ZN(new_n860));
  INV_X1    g0660(.A(new_n439), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n660), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n433), .A2(new_n434), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n427), .A2(new_n439), .ZN(new_n866));
  INV_X1    g0666(.A(new_n660), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n427), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT103), .B1(new_n427), .B2(new_n867), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n864), .B1(new_n870), .B2(KEYINPUT37), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n860), .A2(new_n660), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n436), .B2(new_n442), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n871), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n866), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n863), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n434), .B2(new_n660), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n427), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n428), .B(new_n435), .C1(new_n441), .C2(new_n440), .ZN(new_n889));
  INV_X1    g0689(.A(new_n886), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n880), .A2(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n878), .B(new_n879), .C1(new_n891), .C2(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n876), .A2(new_n877), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n877), .B1(new_n876), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n856), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n809), .B1(new_n807), .B2(new_n817), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n356), .A2(new_n672), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n360), .A2(new_n899), .B1(new_n649), .B2(new_n662), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n871), .A2(new_n873), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n878), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n901), .A2(new_n905), .B1(new_n442), .B2(new_n660), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n725), .A2(new_n728), .A3(new_n449), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n653), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(G330), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT105), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n706), .A2(new_n914), .A3(KEYINPUT31), .A4(new_n662), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n694), .A2(new_n916), .A3(new_n708), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n900), .A2(new_n816), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n878), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT40), .B1(new_n904), .B2(new_n878), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(KEYINPUT40), .B1(new_n923), .B2(new_n920), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n449), .A2(new_n917), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n911), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n910), .B(new_n927), .Z(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n270), .B2(new_n656), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n473), .B1(new_n557), .B2(KEYINPUT35), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n240), .C1(KEYINPUT35), .C2(new_n557), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OAI21_X1  g0732(.A(G77), .B1(new_n224), .B2(new_n228), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n933), .A2(new_n241), .B1(G50), .B2(new_n228), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n655), .A3(new_n293), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n932), .A3(new_n935), .ZN(G367));
  OAI21_X1  g0736(.A(new_n571), .B1(new_n680), .B2(new_n566), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n564), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n564), .A2(new_n679), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n675), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n502), .A2(new_n672), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n632), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n628), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT106), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n941), .B(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n678), .A2(new_n938), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n939), .B1(new_n948), .B2(KEYINPUT42), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n682), .A2(new_n940), .A3(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n951), .B1(KEYINPUT43), .B2(new_n944), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n947), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n685), .B(KEYINPUT41), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n940), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT107), .B1(new_n682), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n678), .A2(new_n958), .A3(new_n681), .A4(new_n940), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n940), .B1(new_n678), .B2(new_n681), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n675), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n673), .A2(new_n674), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n969), .B2(new_n677), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n678), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n671), .A2(KEYINPUT109), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n677), .A2(new_n968), .A3(new_n616), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n675), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n977), .A2(new_n962), .A3(new_n964), .A4(new_n965), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n967), .A2(new_n976), .A3(new_n729), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n955), .B1(new_n979), .B2(new_n729), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n732), .B(KEYINPUT110), .Z(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n953), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n758), .A2(G143), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n738), .A2(G150), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n748), .A2(G68), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G137), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n750), .A2(new_n224), .B1(new_n762), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT113), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n202), .B2(new_n742), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n987), .B(new_n991), .C1(G159), .C2(new_n761), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n302), .C1(new_n217), .C2(new_n753), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n747), .A2(new_n207), .B1(new_n742), .B2(new_n830), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n760), .A2(new_n770), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G311), .C2(new_n758), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT111), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n828), .B2(new_n750), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n739), .A2(G303), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n775), .A2(G97), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n763), .A2(G317), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n793), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT112), .Z(new_n1006));
  OAI21_X1  g0806(.A(new_n993), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n788), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n944), .A2(new_n802), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n792), .B1(new_n211), .B2(new_n363), .C1(new_n251), .C2(new_n796), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1009), .A2(new_n734), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n983), .A2(new_n1012), .ZN(G387));
  INV_X1    g0813(.A(new_n976), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n729), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n685), .B1(new_n976), .B2(new_n729), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n976), .A2(new_n982), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n969), .A2(new_n802), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n779), .A2(new_n202), .B1(new_n762), .B2(new_n277), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n760), .A2(new_n275), .B1(new_n228), .B2(new_n742), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n516), .C2(new_n748), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n793), .B1(G77), .B2(new_n751), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n758), .A2(G159), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1024), .A2(new_n1003), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G322), .A2(new_n758), .B1(new_n761), .B2(G311), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n777), .B2(new_n742), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G317), .B2(new_n739), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT48), .Z(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n830), .B2(new_n747), .C1(new_n770), .C2(new_n750), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT49), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n793), .B1(new_n769), .B2(new_n762), .C1(new_n828), .C2(new_n753), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1027), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n788), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n796), .B1(new_n248), .B2(G45), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n275), .A2(G50), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT50), .Z(new_n1039));
  OAI211_X1 g0839(.A(new_n686), .B(new_n455), .C1(new_n228), .C2(new_n217), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT115), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1037), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n687), .A2(new_n211), .A3(new_n302), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(G107), .B2(new_n211), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n792), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1036), .A2(new_n734), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT117), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1020), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1018), .A2(new_n1019), .A3(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n967), .A2(new_n978), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n685), .A3(new_n979), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n967), .A2(new_n978), .A3(new_n982), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n758), .A2(G317), .B1(G311), .B2(new_n738), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n747), .A2(new_n828), .B1(new_n753), .B2(new_n207), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1058), .A2(new_n302), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n750), .A2(new_n830), .B1(new_n762), .B2(new_n780), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n761), .A2(G303), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1061), .A2(KEYINPUT119), .B1(G294), .B2(new_n743), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n758), .A2(G150), .B1(G159), .B2(new_n738), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n793), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n761), .A2(G50), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n763), .A2(G143), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n747), .A2(new_n217), .B1(new_n742), .B2(new_n275), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n228), .A2(new_n750), .B1(new_n753), .B2(new_n214), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n787), .B1(new_n1065), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n256), .A2(new_n795), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n792), .B(new_n1076), .C1(new_n206), .C2(new_n211), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n735), .B(new_n1075), .C1(KEYINPUT118), .C2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(KEYINPUT118), .B2(new_n1077), .C1(new_n802), .C2(new_n940), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1056), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1055), .A2(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(new_n892), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n879), .B1(new_n904), .B2(new_n878), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT104), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n856), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n897), .B2(new_n900), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n893), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n817), .B1(new_n722), .B2(new_n724), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n810), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n900), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n887), .B1(new_n882), .B2(new_n886), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1092), .A2(new_n1093), .B1(new_n443), .B2(new_n886), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n903), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n856), .B1(new_n1095), .B2(new_n878), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n917), .A2(new_n918), .A3(G330), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n713), .A2(G330), .A3(new_n817), .A4(new_n1090), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1087), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n894), .A2(new_n895), .A3(new_n790), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n760), .A2(new_n207), .B1(new_n206), .B2(new_n742), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n845), .B(new_n331), .C1(new_n214), .C2(new_n750), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n747), .A2(new_n217), .B1(new_n779), .B2(new_n473), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(KEYINPUT120), .B2(new_n1108), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(KEYINPUT120), .B2(new_n1108), .C1(new_n830), .C2(new_n768), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1106), .B(new_n1110), .C1(G294), .C2(new_n763), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n758), .A2(G128), .B1(new_n743), .B2(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n202), .B2(new_n753), .C1(new_n988), .C2(new_n760), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n747), .A2(new_n840), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n751), .A2(G150), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  INV_X1    g0918(.A(G132), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n302), .B1(new_n762), .B2(new_n1118), .C1(new_n779), .C2(new_n1119), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n788), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n851), .A2(new_n275), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n734), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1104), .A2(new_n981), .B1(new_n1105), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n897), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1090), .B1(new_n714), .B2(new_n817), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n1100), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n822), .A2(G330), .A3(new_n917), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n900), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n810), .A3(new_n1088), .A4(new_n1102), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n449), .A2(G330), .A3(new_n917), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n908), .A2(new_n653), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n691), .B1(new_n1104), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1101), .A2(new_n1138), .A3(new_n1103), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1125), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(G378));
  NAND2_X1  g0941(.A1(new_n282), .A2(new_n867), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n320), .B(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n321), .A2(new_n1142), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n320), .B1(new_n282), .B2(new_n867), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n924), .A2(new_n911), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n919), .B1(new_n1095), .B2(new_n878), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT40), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n874), .B2(new_n875), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1153), .A2(new_n1154), .B1(new_n919), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1150), .B1(new_n1156), .B2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n901), .A2(new_n905), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n647), .B2(new_n867), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1085), .B1(new_n1084), .B2(new_n893), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1152), .A2(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n924), .B2(new_n911), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(G330), .A3(new_n1150), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n896), .A4(new_n906), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n981), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1151), .A2(new_n789), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n751), .A2(G77), .B1(new_n763), .B2(G283), .ZN(new_n1167));
  INV_X1    g0967(.A(G41), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n986), .A4(new_n793), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n753), .A2(new_n224), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT121), .Z(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n473), .B2(new_n768), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(G97), .C2(new_n761), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n207), .B2(new_n779), .C1(new_n363), .C2(new_n742), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT58), .Z(new_n1175));
  NOR2_X1   g0975(.A1(G33), .A2(G41), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(G50), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n794), .B2(G41), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n738), .A2(G128), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n760), .B2(new_n1119), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n751), .A2(new_n1112), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n988), .B2(new_n742), .C1(new_n277), .C2(new_n747), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(G125), .C2(new_n758), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT59), .Z(new_n1184));
  INV_X1    g0984(.A(G124), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1176), .B1(new_n762), .B2(new_n1185), .C1(new_n840), .C2(new_n753), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1178), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n788), .B1(new_n1175), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n851), .A2(new_n202), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1166), .A2(new_n734), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT122), .Z(new_n1191));
  NOR2_X1   g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1087), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1099), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1134), .B1(new_n1195), .B2(new_n1138), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT57), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n685), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1139), .A2(new_n1135), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1197), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1192), .B1(new_n1199), .B2(new_n1201), .ZN(G375));
  NOR2_X1   g1002(.A1(new_n768), .A2(new_n1119), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n793), .B(new_n1203), .C1(G137), .C2(new_n739), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n763), .A2(G128), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1171), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G159), .B2(new_n751), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n747), .A2(new_n202), .B1(new_n742), .B2(new_n277), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT124), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n761), .B2(new_n1112), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n762), .A2(new_n777), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n331), .B1(new_n750), .B2(new_n206), .C1(new_n217), .C2(new_n753), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n748), .A2(new_n516), .B1(G283), .B2(new_n738), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1215), .B2(KEYINPUT123), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n761), .A2(new_n468), .B1(G107), .B2(new_n743), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1214), .A2(new_n1218), .B1(new_n758), .B2(G294), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1211), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(new_n788), .B1(new_n228), .B2(new_n851), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n734), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n900), .B2(new_n789), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1132), .B2(new_n982), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n954), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n1138), .ZN(G381));
  OR2_X1    g1027(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1193), .A2(new_n1194), .A3(new_n1136), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1197), .B1(new_n1229), .B2(new_n1134), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n691), .B1(new_n1200), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1228), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1140), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n983), .A2(new_n1012), .A3(new_n1080), .A4(new_n1055), .ZN(new_n1238));
  INV_X1    g1038(.A(G396), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1018), .A2(new_n1239), .A3(new_n1019), .A4(new_n1051), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n1240), .A3(G384), .A4(G381), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(G407));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n661), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G213), .B1(new_n1243), .B2(new_n1236), .ZN(G409));
  AOI22_X1  g1044(.A1(new_n1139), .A2(new_n1135), .B1(new_n1164), .B2(new_n1161), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n954), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1125), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1192), .ZN(new_n1249));
  INV_X1    g1049(.A(G213), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(G343), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1249), .B(new_n1252), .C1(new_n1235), .C2(new_n1140), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT60), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1134), .A2(new_n1128), .A3(KEYINPUT60), .A4(new_n1131), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1136), .A2(new_n1256), .A3(new_n685), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1225), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G384), .B(new_n1225), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1251), .A2(G2897), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1262), .B(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1251), .B1(G375), .B2(G378), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1262), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1249), .A4(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(new_n1266), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(G390), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1238), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1240), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1275), .A2(new_n1272), .A3(KEYINPUT126), .A4(new_n1238), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1271), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1253), .B2(new_n1262), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1279), .A2(KEYINPUT61), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1253), .A2(KEYINPUT125), .A3(new_n1265), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT125), .B1(new_n1253), .B2(new_n1265), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1282), .B(new_n1283), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1249), .A4(new_n1269), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1253), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1269), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1280), .B1(new_n1286), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1200), .A2(new_n1233), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1294), .B(new_n685), .C1(KEYINPUT57), .C2(new_n1245), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1140), .B1(new_n1295), .B2(new_n1192), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1279), .A2(new_n1236), .A3(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1278), .B(new_n1277), .C1(new_n1237), .C2(new_n1296), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1269), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1269), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


