

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799;

  INV_X2 U375 ( .A(G953), .ZN(n790) );
  XNOR2_X1 U376 ( .A(n393), .B(KEYINPUT32), .ZN(n688) );
  NAND2_X2 U377 ( .A1(n663), .A2(n660), .ZN(n659) );
  XNOR2_X2 U378 ( .A(n658), .B(KEYINPUT45), .ZN(n663) );
  XNOR2_X2 U379 ( .A(n662), .B(KEYINPUT87), .ZN(n748) );
  AND2_X2 U380 ( .A1(n618), .A2(n617), .ZN(n662) );
  XNOR2_X2 U381 ( .A(n507), .B(n462), .ZN(n786) );
  XNOR2_X2 U382 ( .A(n537), .B(G134), .ZN(n507) );
  AND2_X1 U383 ( .A1(n644), .A2(n446), .ZN(n445) );
  NOR2_X1 U384 ( .A1(n633), .A2(n365), .ZN(n450) );
  INV_X1 U385 ( .A(n593), .ZN(n717) );
  INV_X1 U386 ( .A(KEYINPUT41), .ZN(n436) );
  NOR2_X1 U387 ( .A1(n422), .A2(n419), .ZN(n610) );
  AND2_X1 U388 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U389 ( .A1(n447), .A2(n445), .ZN(n393) );
  AND2_X1 U390 ( .A1(n452), .A2(n413), .ZN(n373) );
  NAND2_X1 U391 ( .A1(n451), .A2(n450), .ZN(n449) );
  AND2_X1 U392 ( .A1(n725), .A2(n365), .ZN(n415) );
  NAND2_X1 U393 ( .A1(n717), .A2(n716), .ZN(n720) );
  XNOR2_X1 U394 ( .A(n565), .B(KEYINPUT1), .ZN(n572) );
  NOR2_X1 U395 ( .A1(n631), .A2(n728), .ZN(n627) );
  XNOR2_X1 U396 ( .A(n566), .B(n571), .ZN(n619) );
  XNOR2_X1 U397 ( .A(n765), .B(n764), .ZN(n766) );
  XOR2_X1 U398 ( .A(n691), .B(KEYINPUT122), .Z(n692) );
  XNOR2_X1 U399 ( .A(n508), .B(n388), .ZN(n691) );
  XNOR2_X1 U400 ( .A(n456), .B(n530), .ZN(n774) );
  XNOR2_X1 U401 ( .A(n772), .B(KEYINPUT70), .ZN(n536) );
  XNOR2_X1 U402 ( .A(G146), .B(G125), .ZN(n534) );
  XNOR2_X1 U403 ( .A(G104), .B(G107), .ZN(n772) );
  NOR2_X1 U404 ( .A1(n502), .A2(n501), .ZN(n353) );
  NOR2_X1 U405 ( .A1(n502), .A2(n501), .ZN(n552) );
  INV_X1 U406 ( .A(n749), .ZN(n354) );
  NAND2_X2 U407 ( .A1(n410), .A2(n407), .ZN(n565) );
  XNOR2_X2 U408 ( .A(n418), .B(n622), .ZN(n725) );
  INV_X1 U409 ( .A(KEYINPUT86), .ZN(n431) );
  AND2_X1 U410 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U411 ( .A1(n499), .A2(G902), .ZN(n411) );
  NAND2_X1 U412 ( .A1(n421), .A2(n420), .ZN(n419) );
  XNOR2_X1 U413 ( .A(KEYINPUT66), .B(G131), .ZN(n521) );
  NOR2_X1 U414 ( .A1(n748), .A2(n443), .ZN(n440) );
  INV_X1 U415 ( .A(KEYINPUT85), .ZN(n442) );
  NAND2_X1 U416 ( .A1(n691), .A2(n526), .ZN(n511) );
  XNOR2_X1 U417 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n463) );
  INV_X1 U418 ( .A(G119), .ZN(n474) );
  XNOR2_X1 U419 ( .A(n509), .B(n390), .ZN(n389) );
  XNOR2_X1 U420 ( .A(n505), .B(n506), .ZN(n390) );
  INV_X1 U421 ( .A(KEYINPUT7), .ZN(n506) );
  NOR2_X1 U422 ( .A1(n598), .A2(n565), .ZN(n601) );
  XNOR2_X1 U423 ( .A(n592), .B(n366), .ZN(n614) );
  NAND2_X1 U424 ( .A1(n552), .A2(n591), .ZN(n592) );
  XNOR2_X1 U425 ( .A(n416), .B(KEYINPUT110), .ZN(n427) );
  NOR2_X1 U426 ( .A1(n580), .A2(n708), .ZN(n416) );
  NAND2_X1 U427 ( .A1(n379), .A2(n627), .ZN(n378) );
  INV_X1 U428 ( .A(n729), .ZN(n379) );
  BUF_X1 U429 ( .A(n572), .Z(n729) );
  NAND2_X1 U430 ( .A1(n688), .A2(n645), .ZN(n392) );
  INV_X1 U431 ( .A(G237), .ZN(n471) );
  AND2_X1 U432 ( .A1(n355), .A2(n414), .ZN(n413) );
  NAND2_X1 U433 ( .A1(n409), .A2(n526), .ZN(n408) );
  XNOR2_X1 U434 ( .A(G116), .B(G119), .ZN(n466) );
  XOR2_X1 U435 ( .A(KEYINPUT9), .B(KEYINPUT107), .Z(n505) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n516) );
  XNOR2_X1 U437 ( .A(G143), .B(G122), .ZN(n512) );
  XOR2_X1 U438 ( .A(KEYINPUT105), .B(G104), .Z(n513) );
  XOR2_X1 U439 ( .A(KEYINPUT67), .B(G140), .Z(n494) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(G137), .ZN(n461) );
  NAND2_X1 U441 ( .A1(n790), .A2(G224), .ZN(n395) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n544) );
  NOR2_X1 U443 ( .A1(n566), .A2(n581), .ZN(n473) );
  XNOR2_X1 U444 ( .A(n486), .B(n485), .ZN(n577) );
  BUF_X1 U445 ( .A(n748), .Z(n789) );
  XNOR2_X1 U446 ( .A(G137), .B(G128), .ZN(n476) );
  XNOR2_X1 U447 ( .A(KEYINPUT84), .B(KEYINPUT100), .ZN(n475) );
  NAND2_X1 U448 ( .A1(n404), .A2(n441), .ZN(n400) );
  NAND2_X1 U449 ( .A1(n387), .A2(n384), .ZN(n649) );
  NAND2_X1 U450 ( .A1(n385), .A2(KEYINPUT35), .ZN(n384) );
  BUF_X1 U451 ( .A(n566), .Z(n631) );
  XNOR2_X1 U452 ( .A(n504), .B(n389), .ZN(n388) );
  AND2_X1 U453 ( .A1(n668), .A2(G953), .ZN(n771) );
  AND2_X1 U454 ( .A1(n427), .A2(n716), .ZN(n586) );
  INV_X1 U455 ( .A(KEYINPUT42), .ZN(n434) );
  NAND2_X1 U456 ( .A1(n601), .A2(n757), .ZN(n435) );
  INV_X1 U457 ( .A(KEYINPUT40), .ZN(n437) );
  INV_X1 U458 ( .A(KEYINPUT36), .ZN(n455) );
  NAND2_X1 U459 ( .A1(n377), .A2(n376), .ZN(n629) );
  INV_X1 U460 ( .A(n378), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n624), .B(KEYINPUT77), .ZN(n355) );
  XOR2_X1 U462 ( .A(n530), .B(n468), .Z(n356) );
  XOR2_X1 U463 ( .A(n477), .B(n476), .Z(n357) );
  AND2_X1 U464 ( .A1(n487), .A2(G217), .ZN(n358) );
  XNOR2_X1 U465 ( .A(n428), .B(KEYINPUT75), .ZN(n753) );
  AND2_X1 U466 ( .A1(n430), .A2(G472), .ZN(n359) );
  AND2_X1 U467 ( .A1(n430), .A2(G475), .ZN(n360) );
  AND2_X1 U468 ( .A1(n430), .A2(G210), .ZN(n361) );
  NAND2_X1 U469 ( .A1(n605), .A2(n604), .ZN(n362) );
  AND2_X1 U470 ( .A1(n631), .A2(n630), .ZN(n363) );
  AND2_X1 U471 ( .A1(n585), .A2(n716), .ZN(n364) );
  XOR2_X1 U472 ( .A(KEYINPUT73), .B(KEYINPUT34), .Z(n365) );
  XNOR2_X1 U473 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n366) );
  XOR2_X1 U474 ( .A(n553), .B(KEYINPUT19), .Z(n367) );
  INV_X1 U475 ( .A(KEYINPUT35), .ZN(n414) );
  AND2_X1 U476 ( .A1(n441), .A2(KEYINPUT64), .ZN(n368) );
  INV_X1 U477 ( .A(KEYINPUT64), .ZN(n444) );
  BUF_X1 U478 ( .A(n725), .Z(n369) );
  INV_X1 U479 ( .A(n460), .ZN(n446) );
  XNOR2_X1 U480 ( .A(n370), .B(n564), .ZN(n569) );
  NOR2_X1 U481 ( .A1(n623), .A2(n562), .ZN(n370) );
  NAND2_X1 U482 ( .A1(n401), .A2(n400), .ZN(n402) );
  AND2_X1 U483 ( .A1(n405), .A2(n444), .ZN(n401) );
  AND2_X1 U484 ( .A1(n452), .A2(n355), .ZN(n386) );
  BUF_X1 U485 ( .A(n665), .Z(n371) );
  XNOR2_X1 U486 ( .A(n538), .B(n395), .ZN(n394) );
  XNOR2_X1 U487 ( .A(G104), .B(G107), .ZN(n372) );
  XNOR2_X1 U488 ( .A(n786), .B(G146), .ZN(n374) );
  XNOR2_X1 U489 ( .A(n786), .B(G146), .ZN(n497) );
  XNOR2_X1 U490 ( .A(n532), .B(n529), .ZN(n456) );
  XNOR2_X1 U491 ( .A(n535), .B(n536), .ZN(n458) );
  INV_X1 U492 ( .A(n454), .ZN(n375) );
  INV_X1 U493 ( .A(n454), .ZN(n439) );
  NAND2_X1 U494 ( .A1(n406), .A2(n430), .ZN(n454) );
  INV_X1 U495 ( .A(n633), .ZN(n377) );
  NAND2_X1 U496 ( .A1(n739), .A2(n378), .ZN(n740) );
  NAND2_X1 U497 ( .A1(n381), .A2(n380), .ZN(n383) );
  INV_X1 U498 ( .A(n415), .ZN(n380) );
  NAND2_X1 U499 ( .A1(n449), .A2(n373), .ZN(n381) );
  NAND2_X1 U500 ( .A1(n383), .A2(n382), .ZN(n387) );
  NAND2_X1 U501 ( .A1(n415), .A2(n414), .ZN(n382) );
  NAND2_X1 U502 ( .A1(n449), .A2(n386), .ZN(n385) );
  INV_X1 U503 ( .A(n725), .ZN(n451) );
  BUF_X2 U504 ( .A(n588), .Z(n583) );
  NAND2_X1 U505 ( .A1(n391), .A2(n432), .ZN(n405) );
  NAND2_X1 U506 ( .A1(n440), .A2(n391), .ZN(n404) );
  XNOR2_X2 U507 ( .A(n659), .B(n431), .ZN(n391) );
  XNOR2_X2 U508 ( .A(n392), .B(KEYINPUT93), .ZN(n653) );
  XNOR2_X1 U509 ( .A(n537), .B(n394), .ZN(n459) );
  XNOR2_X2 U510 ( .A(n396), .B(G128), .ZN(n537) );
  XNOR2_X2 U511 ( .A(G143), .B(KEYINPUT78), .ZN(n396) );
  AND2_X2 U512 ( .A1(n398), .A2(n397), .ZN(n403) );
  NAND2_X1 U513 ( .A1(n404), .A2(n368), .ZN(n397) );
  NAND2_X1 U514 ( .A1(n399), .A2(KEYINPUT64), .ZN(n398) );
  INV_X1 U515 ( .A(n405), .ZN(n399) );
  NAND2_X2 U516 ( .A1(n403), .A2(n402), .ZN(n406) );
  NAND2_X1 U517 ( .A1(n406), .A2(n359), .ZN(n667) );
  NAND2_X1 U518 ( .A1(n406), .A2(n360), .ZN(n674) );
  NAND2_X1 U519 ( .A1(n406), .A2(n361), .ZN(n683) );
  OR2_X1 U520 ( .A1(n762), .A2(n408), .ZN(n407) );
  INV_X1 U521 ( .A(n499), .ZN(n409) );
  NAND2_X1 U522 ( .A1(n762), .A2(n499), .ZN(n412) );
  INV_X1 U523 ( .A(n572), .ZN(n620) );
  XNOR2_X1 U524 ( .A(n767), .B(n766), .ZN(n417) );
  XNOR2_X1 U525 ( .A(n497), .B(n356), .ZN(n665) );
  NAND2_X1 U526 ( .A1(n621), .A2(n620), .ZN(n418) );
  NOR2_X1 U527 ( .A1(n417), .A2(n771), .ZN(G54) );
  NAND2_X1 U528 ( .A1(n363), .A2(n500), .ZN(n632) );
  INV_X1 U529 ( .A(n565), .ZN(n500) );
  INV_X1 U530 ( .A(n797), .ZN(n424) );
  XNOR2_X2 U531 ( .A(n438), .B(n437), .ZN(n797) );
  XNOR2_X2 U532 ( .A(n435), .B(n434), .ZN(n799) );
  NAND2_X1 U533 ( .A1(n797), .A2(KEYINPUT46), .ZN(n420) );
  NAND2_X1 U534 ( .A1(n799), .A2(KEYINPUT46), .ZN(n421) );
  NAND2_X1 U535 ( .A1(n362), .A2(n423), .ZN(n422) );
  NAND2_X1 U536 ( .A1(n425), .A2(n424), .ZN(n423) );
  NOR2_X1 U537 ( .A1(n799), .A2(KEYINPUT46), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n427), .A2(n364), .ZN(n426) );
  XNOR2_X1 U539 ( .A(n426), .B(n455), .ZN(n587) );
  NAND2_X1 U540 ( .A1(n429), .A2(n354), .ZN(n428) );
  AND2_X1 U541 ( .A1(n662), .A2(KEYINPUT2), .ZN(n429) );
  INV_X1 U542 ( .A(n753), .ZN(n430) );
  NOR2_X1 U543 ( .A1(n748), .A2(KEYINPUT85), .ZN(n432) );
  XNOR2_X2 U544 ( .A(n583), .B(n589), .ZN(n593) );
  XNOR2_X2 U545 ( .A(n433), .B(n543), .ZN(n588) );
  OR2_X2 U546 ( .A1(n681), .A2(n660), .ZN(n433) );
  NAND2_X1 U547 ( .A1(n614), .A2(n704), .ZN(n438) );
  XNOR2_X2 U548 ( .A(n594), .B(n436), .ZN(n757) );
  NAND2_X1 U549 ( .A1(n375), .A2(G469), .ZN(n767) );
  NAND2_X1 U550 ( .A1(n439), .A2(G478), .ZN(n693) );
  NAND2_X1 U551 ( .A1(n661), .A2(n442), .ZN(n441) );
  INV_X1 U552 ( .A(n661), .ZN(n443) );
  NOR2_X1 U553 ( .A1(n569), .A2(n460), .ZN(n448) );
  INV_X1 U554 ( .A(n569), .ZN(n447) );
  NAND2_X1 U555 ( .A1(n448), .A2(n729), .ZN(n573) );
  NAND2_X1 U556 ( .A1(n633), .A2(n365), .ZN(n452) );
  XNOR2_X2 U557 ( .A(n470), .B(n469), .ZN(n566) );
  NOR2_X1 U558 ( .A1(n454), .A2(n453), .ZN(n769) );
  INV_X1 U559 ( .A(G217), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n457), .B(n774), .ZN(n681) );
  XNOR2_X1 U561 ( .A(n459), .B(n458), .ZN(n457) );
  INV_X1 U562 ( .A(n619), .ZN(n460) );
  BUF_X1 U563 ( .A(n649), .Z(n690) );
  NOR2_X1 U564 ( .A1(n665), .A2(G902), .ZN(n470) );
  BUF_X1 U565 ( .A(n577), .Z(n731) );
  XNOR2_X1 U566 ( .A(n521), .B(n461), .ZN(n462) );
  XNOR2_X1 U567 ( .A(G101), .B(G113), .ZN(n464) );
  XNOR2_X1 U568 ( .A(n464), .B(n463), .ZN(n530) );
  NOR2_X1 U569 ( .A1(G953), .A2(G237), .ZN(n514) );
  NAND2_X1 U570 ( .A1(n514), .A2(G210), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n465), .B(KEYINPUT5), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U573 ( .A(G472), .B(KEYINPUT103), .Z(n469) );
  INV_X1 U574 ( .A(G902), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n526), .A2(n471), .ZN(n540) );
  AND2_X1 U576 ( .A1(n540), .A2(G214), .ZN(n581) );
  XNOR2_X1 U577 ( .A(KEYINPUT30), .B(KEYINPUT111), .ZN(n472) );
  XNOR2_X1 U578 ( .A(n473), .B(n472), .ZN(n502) );
  XNOR2_X1 U579 ( .A(n474), .B(G110), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(n475), .ZN(n478) );
  XOR2_X1 U581 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n477) );
  XNOR2_X1 U582 ( .A(n478), .B(n357), .ZN(n481) );
  NAND2_X1 U583 ( .A1(G234), .A2(n790), .ZN(n479) );
  XOR2_X1 U584 ( .A(KEYINPUT8), .B(n479), .Z(n503) );
  NAND2_X1 U585 ( .A1(G221), .A2(n503), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT10), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n494), .B(n523), .ZN(n787) );
  XNOR2_X1 U589 ( .A(n482), .B(n787), .ZN(n768) );
  NAND2_X1 U590 ( .A1(n768), .A2(n526), .ZN(n486) );
  XOR2_X1 U591 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n484) );
  XNOR2_X1 U592 ( .A(G902), .B(KEYINPUT15), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n539), .A2(G234), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n483), .B(KEYINPUT20), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n484), .B(n358), .ZN(n485) );
  AND2_X1 U596 ( .A1(n487), .A2(G221), .ZN(n489) );
  XNOR2_X1 U597 ( .A(KEYINPUT102), .B(KEYINPUT21), .ZN(n488) );
  XNOR2_X1 U598 ( .A(n489), .B(n488), .ZN(n732) );
  NAND2_X1 U599 ( .A1(n577), .A2(n732), .ZN(n728) );
  INV_X1 U600 ( .A(n728), .ZN(n630) );
  XNOR2_X1 U601 ( .A(G101), .B(G110), .ZN(n490) );
  XNOR2_X1 U602 ( .A(KEYINPUT99), .B(n490), .ZN(n492) );
  NAND2_X1 U603 ( .A1(n790), .A2(G227), .ZN(n491) );
  XNOR2_X1 U604 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U606 ( .A(n495), .B(n536), .ZN(n496) );
  XNOR2_X1 U607 ( .A(n374), .B(n496), .ZN(n762) );
  INV_X1 U608 ( .A(KEYINPUT68), .ZN(n498) );
  XNOR2_X1 U609 ( .A(n498), .B(G469), .ZN(n499) );
  NAND2_X1 U610 ( .A1(n630), .A2(n500), .ZN(n501) );
  NAND2_X1 U611 ( .A1(G217), .A2(n503), .ZN(n504) );
  BUF_X1 U612 ( .A(n507), .Z(n508) );
  XNOR2_X2 U613 ( .A(G122), .B(G116), .ZN(n531) );
  XNOR2_X1 U614 ( .A(n531), .B(G107), .ZN(n509) );
  XNOR2_X1 U615 ( .A(KEYINPUT108), .B(G478), .ZN(n510) );
  XNOR2_X1 U616 ( .A(n511), .B(n510), .ZN(n576) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n518) );
  NAND2_X1 U618 ( .A1(G214), .A2(n514), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n525) );
  INV_X1 U621 ( .A(G113), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n519), .B(G140), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U625 ( .A(n525), .B(n524), .ZN(n672) );
  NAND2_X1 U626 ( .A1(n672), .A2(n526), .ZN(n528) );
  XOR2_X1 U627 ( .A(KEYINPUT13), .B(G475), .Z(n527) );
  XNOR2_X1 U628 ( .A(n528), .B(n527), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n576), .A2(n575), .ZN(n624) );
  XNOR2_X1 U630 ( .A(n531), .B(KEYINPUT16), .ZN(n532) );
  XNOR2_X1 U631 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n533) );
  XNOR2_X1 U632 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U633 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n538) );
  INV_X1 U634 ( .A(n539), .ZN(n660) );
  NAND2_X1 U635 ( .A1(n540), .A2(G210), .ZN(n542) );
  INV_X1 U636 ( .A(KEYINPUT79), .ZN(n541) );
  XNOR2_X1 U637 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U638 ( .A(n583), .ZN(n585) );
  XNOR2_X1 U639 ( .A(n544), .B(KEYINPUT96), .ZN(n545) );
  XNOR2_X1 U640 ( .A(KEYINPUT14), .B(n545), .ZN(n546) );
  NAND2_X1 U641 ( .A1(G952), .A2(n546), .ZN(n747) );
  NOR2_X1 U642 ( .A1(G953), .A2(n747), .ZN(n557) );
  NAND2_X1 U643 ( .A1(G902), .A2(n546), .ZN(n555) );
  OR2_X1 U644 ( .A1(n790), .A2(n555), .ZN(n547) );
  NOR2_X1 U645 ( .A1(G900), .A2(n547), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n557), .A2(n548), .ZN(n590) );
  INV_X1 U647 ( .A(n590), .ZN(n549) );
  NAND2_X1 U648 ( .A1(n585), .A2(n549), .ZN(n550) );
  NOR2_X1 U649 ( .A1(n624), .A2(n550), .ZN(n551) );
  NAND2_X1 U650 ( .A1(n353), .A2(n551), .ZN(n607) );
  XNOR2_X1 U651 ( .A(n607), .B(G143), .ZN(G45) );
  NOR2_X2 U652 ( .A1(n588), .A2(n581), .ZN(n554) );
  INV_X1 U653 ( .A(KEYINPUT65), .ZN(n553) );
  XNOR2_X1 U654 ( .A(n554), .B(n367), .ZN(n599) );
  XNOR2_X1 U655 ( .A(G898), .B(KEYINPUT97), .ZN(n780) );
  NAND2_X1 U656 ( .A1(G953), .A2(n780), .ZN(n775) );
  NOR2_X1 U657 ( .A1(n555), .A2(n775), .ZN(n556) );
  OR2_X1 U658 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n558), .B(KEYINPUT98), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n599), .A2(n559), .ZN(n560) );
  XNOR2_X1 U661 ( .A(n560), .B(KEYINPUT0), .ZN(n623) );
  OR2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n719) );
  INV_X1 U663 ( .A(n719), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n561), .A2(n732), .ZN(n562) );
  INV_X1 U665 ( .A(KEYINPUT74), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n563), .B(KEYINPUT22), .ZN(n564) );
  INV_X1 U667 ( .A(n631), .ZN(n734) );
  OR2_X1 U668 ( .A1(n734), .A2(n731), .ZN(n567) );
  OR2_X1 U669 ( .A1(n620), .A2(n567), .ZN(n568) );
  OR2_X1 U670 ( .A1(n569), .A2(n568), .ZN(n645) );
  XNOR2_X1 U671 ( .A(G110), .B(KEYINPUT114), .ZN(n570) );
  XNOR2_X1 U672 ( .A(n645), .B(n570), .ZN(G12) );
  INV_X1 U673 ( .A(KEYINPUT6), .ZN(n571) );
  XNOR2_X1 U674 ( .A(n573), .B(KEYINPUT89), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n574), .A2(n731), .ZN(n637) );
  XNOR2_X1 U676 ( .A(n637), .B(G101), .ZN(G3) );
  XNOR2_X1 U677 ( .A(n575), .B(KEYINPUT106), .ZN(n603) );
  INV_X1 U678 ( .A(n576), .ZN(n602) );
  AND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n704) );
  INV_X1 U680 ( .A(n704), .ZN(n708) );
  NOR2_X1 U681 ( .A1(n590), .A2(n577), .ZN(n578) );
  NAND2_X1 U682 ( .A1(n732), .A2(n578), .ZN(n595) );
  NOR2_X1 U683 ( .A1(n619), .A2(n595), .ZN(n579) );
  XNOR2_X1 U684 ( .A(n579), .B(KEYINPUT109), .ZN(n580) );
  INV_X1 U685 ( .A(n581), .ZN(n716) );
  NAND2_X1 U686 ( .A1(n586), .A2(n729), .ZN(n582) );
  XNOR2_X1 U687 ( .A(n582), .B(KEYINPUT43), .ZN(n584) );
  NAND2_X1 U688 ( .A1(n584), .A2(n583), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(G140), .ZN(G42) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT94), .ZN(n643) );
  AND2_X1 U691 ( .A1(n587), .A2(n643), .ZN(n713) );
  XNOR2_X1 U692 ( .A(n713), .B(KEYINPUT88), .ZN(n612) );
  INV_X1 U693 ( .A(KEYINPUT38), .ZN(n589) );
  NOR2_X1 U694 ( .A1(n593), .A2(n590), .ZN(n591) );
  NOR2_X2 U695 ( .A1(n719), .A2(n720), .ZN(n594) );
  NOR2_X1 U696 ( .A1(n631), .A2(n595), .ZN(n597) );
  XOR2_X1 U697 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n596) );
  XNOR2_X1 U698 ( .A(n597), .B(n596), .ZN(n598) );
  BUF_X1 U699 ( .A(n599), .Z(n600) );
  NAND2_X1 U700 ( .A1(n601), .A2(n600), .ZN(n700) );
  XNOR2_X1 U701 ( .A(n700), .B(KEYINPUT47), .ZN(n605) );
  NOR2_X1 U702 ( .A1(n603), .A2(n602), .ZN(n701) );
  NOR2_X1 U703 ( .A1(n704), .A2(n701), .ZN(n721) );
  XNOR2_X1 U704 ( .A(KEYINPUT83), .B(n721), .ZN(n634) );
  OR2_X1 U705 ( .A1(n700), .A2(n634), .ZN(n604) );
  NAND2_X1 U706 ( .A1(n721), .A2(KEYINPUT47), .ZN(n606) );
  NAND2_X1 U707 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U708 ( .A(n608), .B(KEYINPUT80), .Z(n609) );
  NAND2_X1 U709 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X2 U710 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U711 ( .A(n613), .B(KEYINPUT48), .ZN(n618) );
  AND2_X1 U712 ( .A1(n614), .A2(n701), .ZN(n715) );
  INV_X1 U713 ( .A(n715), .ZN(n615) );
  AND2_X1 U714 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U715 ( .A1(n619), .A2(n728), .ZN(n621) );
  XNOR2_X1 U716 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n622) );
  BUF_X2 U717 ( .A(n623), .Z(n633) );
  NAND2_X1 U718 ( .A1(n649), .A2(KEYINPUT44), .ZN(n626) );
  INV_X1 U719 ( .A(KEYINPUT91), .ZN(n625) );
  XNOR2_X1 U720 ( .A(n626), .B(n625), .ZN(n639) );
  XOR2_X1 U721 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n628) );
  XNOR2_X1 U722 ( .A(n629), .B(n628), .ZN(n711) );
  OR2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n696) );
  NAND2_X1 U724 ( .A1(n711), .A2(n696), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n641) );
  INV_X1 U727 ( .A(KEYINPUT90), .ZN(n640) );
  XNOR2_X1 U728 ( .A(n641), .B(n640), .ZN(n657) );
  INV_X1 U729 ( .A(n731), .ZN(n642) );
  AND2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n644) );
  INV_X1 U731 ( .A(n653), .ZN(n648) );
  OR2_X1 U732 ( .A1(n649), .A2(KEYINPUT92), .ZN(n646) );
  INV_X1 U733 ( .A(KEYINPUT44), .ZN(n650) );
  AND2_X1 U734 ( .A1(n646), .A2(n650), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n650), .A2(KEYINPUT92), .ZN(n651) );
  OR2_X1 U737 ( .A1(n690), .A2(n651), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n660), .A2(KEYINPUT2), .ZN(n661) );
  XNOR2_X1 U742 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n371), .B(n664), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n667), .B(n666), .ZN(n669) );
  INV_X1 U745 ( .A(G952), .ZN(n668) );
  INV_X1 U746 ( .A(n771), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n669), .A2(n684), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U749 ( .A(KEYINPUT95), .B(KEYINPUT59), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n675), .A2(n684), .ZN(n677) );
  INV_X1 U753 ( .A(KEYINPUT60), .ZN(n676) );
  XNOR2_X1 U754 ( .A(n677), .B(n676), .ZN(G60) );
  XOR2_X1 U755 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n679) );
  XNOR2_X1 U756 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U760 ( .A1(n685), .A2(n684), .ZN(n687) );
  INV_X1 U761 ( .A(KEYINPUT56), .ZN(n686) );
  XNOR2_X1 U762 ( .A(n687), .B(n686), .ZN(G51) );
  BUF_X1 U763 ( .A(n688), .Z(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(G119), .ZN(G21) );
  XOR2_X1 U765 ( .A(n690), .B(G122), .Z(G24) );
  XNOR2_X1 U766 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U767 ( .A1(n694), .A2(n771), .ZN(G63) );
  NOR2_X1 U768 ( .A1(n708), .A2(n696), .ZN(n695) );
  XOR2_X1 U769 ( .A(G104), .B(n695), .Z(G6) );
  INV_X1 U770 ( .A(n701), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n710), .A2(n696), .ZN(n698) );
  XNOR2_X1 U772 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n697) );
  XNOR2_X1 U773 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U774 ( .A(G107), .B(n699), .ZN(G9) );
  XOR2_X1 U775 ( .A(G128), .B(KEYINPUT29), .Z(n703) );
  INV_X1 U776 ( .A(n700), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n705), .A2(n701), .ZN(n702) );
  XNOR2_X1 U778 ( .A(n703), .B(n702), .ZN(G30) );
  XOR2_X1 U779 ( .A(G146), .B(KEYINPUT115), .Z(n707) );
  NAND2_X1 U780 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U781 ( .A(n707), .B(n706), .ZN(G48) );
  NOR2_X1 U782 ( .A1(n711), .A2(n708), .ZN(n709) );
  XOR2_X1 U783 ( .A(G113), .B(n709), .Z(G15) );
  NOR2_X1 U784 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U785 ( .A(G116), .B(n712), .Z(G18) );
  XNOR2_X1 U786 ( .A(G125), .B(n713), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n714), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U788 ( .A(G134), .B(n715), .Z(G36) );
  NOR2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U793 ( .A(KEYINPUT118), .B(n724), .Z(n726) );
  INV_X1 U794 ( .A(n369), .ZN(n756) );
  NAND2_X1 U795 ( .A1(n726), .A2(n756), .ZN(n727) );
  XNOR2_X1 U796 ( .A(n727), .B(KEYINPUT119), .ZN(n744) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U798 ( .A(n730), .B(KEYINPUT50), .ZN(n738) );
  NOR2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U800 ( .A(KEYINPUT49), .B(n733), .Z(n735) );
  NOR2_X1 U801 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U802 ( .A(n736), .B(KEYINPUT116), .ZN(n737) );
  NAND2_X1 U803 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U804 ( .A(KEYINPUT51), .B(n740), .Z(n741) );
  NAND2_X1 U805 ( .A1(n757), .A2(n741), .ZN(n742) );
  XNOR2_X1 U806 ( .A(KEYINPUT117), .B(n742), .ZN(n743) );
  NOR2_X1 U807 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U808 ( .A(n745), .B(KEYINPUT52), .ZN(n746) );
  NOR2_X1 U809 ( .A1(n747), .A2(n746), .ZN(n755) );
  INV_X1 U810 ( .A(n663), .ZN(n749) );
  OR2_X1 U811 ( .A1(n789), .A2(n749), .ZN(n751) );
  XOR2_X1 U812 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n750) );
  AND2_X1 U813 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U814 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U815 ( .A1(n755), .A2(n754), .ZN(n759) );
  NAND2_X1 U816 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U817 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U818 ( .A1(n760), .A2(G953), .ZN(n761) );
  XNOR2_X1 U819 ( .A(n761), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U820 ( .A(n762), .Z(n765) );
  XNOR2_X1 U821 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n763) );
  XNOR2_X1 U822 ( .A(n763), .B(KEYINPUT57), .ZN(n764) );
  XNOR2_X1 U823 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U824 ( .A1(n770), .A2(n771), .ZN(G66) );
  XNOR2_X1 U825 ( .A(n372), .B(KEYINPUT125), .ZN(n773) );
  XNOR2_X1 U826 ( .A(n774), .B(n773), .ZN(n776) );
  NAND2_X1 U827 ( .A1(n776), .A2(n775), .ZN(n785) );
  NAND2_X1 U828 ( .A1(G224), .A2(G953), .ZN(n777) );
  XNOR2_X1 U829 ( .A(n777), .B(KEYINPUT123), .ZN(n778) );
  XNOR2_X1 U830 ( .A(n778), .B(KEYINPUT61), .ZN(n779) );
  NOR2_X1 U831 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U832 ( .A1(n354), .A2(n790), .ZN(n781) );
  XOR2_X1 U833 ( .A(KEYINPUT124), .B(n781), .Z(n782) );
  NOR2_X1 U834 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U835 ( .A(n785), .B(n784), .ZN(G69) );
  XNOR2_X1 U836 ( .A(n787), .B(KEYINPUT126), .ZN(n788) );
  XOR2_X1 U837 ( .A(n786), .B(n788), .Z(n792) );
  XNOR2_X1 U838 ( .A(n792), .B(n789), .ZN(n791) );
  NAND2_X1 U839 ( .A1(n791), .A2(n790), .ZN(n796) );
  XNOR2_X1 U840 ( .A(G227), .B(n792), .ZN(n793) );
  NAND2_X1 U841 ( .A1(n793), .A2(G900), .ZN(n794) );
  NAND2_X1 U842 ( .A1(G953), .A2(n794), .ZN(n795) );
  NAND2_X1 U843 ( .A1(n796), .A2(n795), .ZN(G72) );
  XNOR2_X1 U844 ( .A(G131), .B(KEYINPUT127), .ZN(n798) );
  XNOR2_X1 U845 ( .A(n798), .B(n797), .ZN(G33) );
  XOR2_X1 U846 ( .A(G137), .B(n799), .Z(G39) );
endmodule

