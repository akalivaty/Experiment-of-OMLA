//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n210), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n212), .A2(KEYINPUT28), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT28), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n209), .B(new_n211), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  OAI211_X1 g018(.A(KEYINPUT25), .B(new_n217), .C1(new_n219), .C2(new_n210), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n221), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n218), .A2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(new_n204), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n206), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n228), .A2(new_n231), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G169gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n216), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G134gat), .ZN(new_n251));
  INV_X1    g050(.A(G134gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(G127gat), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n249), .A2(KEYINPUT1), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n254), .A2(new_n262), .A3(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n226), .A2(new_n244), .A3(new_n245), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n229), .B1(new_n271), .B2(new_n241), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n225), .A3(new_n235), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n267), .A2(new_n273), .A3(new_n216), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n270), .A4(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n203), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT33), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G43gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT69), .ZN(new_n282));
  XOR2_X1   g081(.A(G71gat), .B(G99gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT34), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI221_X4 g088(.A(new_n203), .B1(KEYINPUT33), .B2(new_n284), .C1(new_n277), .C2(new_n278), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n277), .A2(new_n278), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n284), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n285), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n288), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n269), .A2(new_n274), .ZN(new_n299));
  OAI22_X1  g098(.A1(new_n299), .A2(new_n270), .B1(new_n287), .B2(KEYINPUT34), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n291), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n289), .B1(new_n286), .B2(new_n290), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n296), .A2(new_n288), .A3(new_n297), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n202), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT71), .B(G211gat), .Z(new_n308));
  INV_X1    g107(.A(G218gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n312), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G141gat), .B(G148gat), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n318), .B(new_n321), .C1(new_n322), .C2(KEYINPUT2), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n318), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n323), .A2(new_n324), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT3), .B1(new_n316), .B2(new_n334), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n323), .A2(new_n332), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G22gat), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT31), .B(G50gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  AOI22_X1  g146(.A1(new_n340), .A2(new_n342), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n344), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT79), .Z(new_n350));
  AND3_X1   g149(.A1(new_n343), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n343), .B2(new_n348), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n273), .A2(new_n216), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n334), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n273), .B2(new_n216), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n317), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n248), .A2(new_n360), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n273), .A2(new_n216), .A3(new_n358), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n316), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n366), .A3(KEYINPUT73), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .A4(new_n316), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n357), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n369), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n357), .B(KEYINPUT74), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI22_X1  g172(.A1(new_n370), .A2(KEYINPUT30), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n370), .A2(KEYINPUT30), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n323), .A2(new_n254), .A3(new_n332), .A4(new_n262), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n265), .A2(new_n339), .A3(new_n266), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(new_n382), .C1(KEYINPUT4), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n263), .A3(new_n333), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n392));
  AND4_X1   g191(.A1(new_n323), .A2(new_n254), .A3(new_n332), .A4(new_n262), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n378), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(KEYINPUT4), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n338), .A2(new_n263), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n388), .B1(new_n400), .B2(new_n378), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT76), .B1(new_n401), .B2(new_n385), .ZN(new_n402));
  INV_X1    g201(.A(new_n388), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n323), .A2(new_n332), .B1(new_n254), .B2(new_n262), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n393), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n390), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n390), .B(new_n416), .C1(new_n399), .C2(new_n408), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n354), .B1(new_n377), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n300), .B1(new_n291), .B2(new_n298), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n303), .A2(new_n302), .A3(new_n304), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n306), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n388), .B1(new_n384), .B2(new_n387), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n378), .A3(new_n388), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT39), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n413), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(KEYINPUT40), .A3(new_n433), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n414), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n353), .B1(new_n376), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT38), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n367), .A2(KEYINPUT37), .A3(new_n369), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(new_n357), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n371), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n418), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n372), .A2(new_n440), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n363), .A2(new_n366), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n370), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n414), .A2(KEYINPUT80), .A3(new_n415), .A4(new_n417), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n447), .A2(new_n451), .A3(new_n419), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n453), .B2(KEYINPUT81), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n419), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n447), .A4(new_n451), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n427), .B(new_n439), .C1(new_n454), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(KEYINPUT81), .ZN(new_n459));
  INV_X1    g258(.A(new_n445), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n439), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT82), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n426), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n354), .B1(new_n423), .B2(new_n424), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n377), .A2(new_n421), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n468), .B(new_n377), .C1(new_n447), .C2(new_n455), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n467), .A2(KEYINPUT35), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT84), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n306), .A2(new_n425), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n427), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n461), .A2(KEYINPUT82), .A3(new_n462), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n422), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n465), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G8gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT16), .ZN(new_n487));
  AOI21_X1  g286(.A(G1gat), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n486), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G43gat), .B(G50gat), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n494), .A2(KEYINPUT87), .A3(KEYINPUT15), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT15), .B1(new_n494), .B2(KEYINPUT87), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n493), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(KEYINPUT17), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n493), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT89), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n491), .A2(new_n492), .ZN(new_n517));
  INV_X1    g316(.A(new_n513), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n504), .B2(new_n506), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n493), .A2(new_n507), .B1(G229gat), .B2(G233gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT90), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n509), .B(KEYINPUT13), .Z(new_n526));
  INV_X1    g325(.A(new_n508), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n493), .A2(new_n507), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(new_n522), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n516), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT91), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n523), .A3(new_n533), .A4(new_n516), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n529), .B(new_n535), .C1(new_n530), .C2(new_n516), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n525), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549));
  INV_X1    g348(.A(new_n524), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n529), .B(new_n544), .C1(new_n530), .C2(new_n516), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .A3(new_n524), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n545), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n564), .B2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n563), .A2(new_n566), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n573), .A2(new_n561), .A3(new_n567), .A4(new_n569), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G71gat), .B(G78gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n577), .A3(new_n578), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n560), .B1(new_n575), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n583), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n572), .A3(new_n574), .A4(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n567), .A3(new_n569), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n562), .A2(KEYINPUT99), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  XOR2_X1   g391(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n584), .B(KEYINPUT94), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n559), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n558), .B1(new_n588), .B2(new_n592), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n598), .B2(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G127gat), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n493), .B1(new_n596), .B2(KEYINPUT21), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n575), .B2(new_n507), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n518), .A2(new_n519), .ZN(new_n626));
  OAI22_X1  g425(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n575), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  AND3_X1   g433(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n629), .B2(new_n630), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n482), .A2(new_n557), .A3(new_n607), .A4(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n421), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g441(.A(new_n489), .B1(new_n640), .B2(new_n377), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n639), .A2(new_n376), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  OAI21_X1  g446(.A(G15gat), .B1(new_n639), .B2(new_n472), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n301), .A2(new_n305), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n639), .B2(new_n650), .ZN(G1326gat));
  OAI21_X1  g450(.A(KEYINPUT101), .B1(new_n639), .B2(new_n353), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n639), .A2(KEYINPUT101), .A3(new_n353), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT102), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n652), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n655), .B2(new_n658), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n637), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n471), .B2(new_n481), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n620), .A2(new_n606), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n548), .A2(new_n555), .A3(new_n556), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(G29gat), .A3(new_n420), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT45), .Z(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(new_n476), .B2(new_n479), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n664), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n668), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(KEYINPUT103), .A3(new_n668), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n678), .A2(new_n421), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n671), .B1(new_n680), .B2(new_n496), .ZN(G1328gat));
  NOR3_X1   g480(.A1(new_n669), .A2(G36gat), .A3(new_n376), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n678), .A2(new_n377), .A3(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n497), .ZN(G1329gat));
  INV_X1    g484(.A(new_n649), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n666), .A2(G43gat), .A3(new_n663), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n482), .A2(new_n686), .A3(new_n557), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n472), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n678), .A2(new_n690), .A3(new_n679), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n691), .B2(G43gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(KEYINPUT47), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n690), .A3(new_n668), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G43gat), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n697));
  OAI22_X1  g496(.A1(new_n692), .A2(KEYINPUT47), .B1(new_n696), .B2(new_n697), .ZN(G1330gat));
  NOR3_X1   g497(.A1(new_n669), .A2(G50gat), .A3(new_n353), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT48), .B(G50gat), .C1(new_n676), .C2(new_n353), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n678), .A2(new_n354), .A3(new_n679), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(G50gat), .B1(new_n700), .B2(new_n699), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g506(.A1(new_n638), .A2(new_n667), .A3(new_n606), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT106), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n479), .B2(new_n476), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n421), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n376), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(G1333gat));
  NAND3_X1  g516(.A1(new_n710), .A2(G71gat), .A3(new_n690), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n649), .B(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n721), .B2(G71gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g522(.A1(new_n710), .A2(new_n354), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n621), .A2(new_n667), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n637), .B(new_n727), .C1(new_n464), .C2(new_n470), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT109), .B1(new_n729), .B2(KEYINPUT51), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n672), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n727), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n607), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n564), .A3(new_n421), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n726), .A2(new_n607), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n675), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n421), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n564), .ZN(G1336gat));
  AOI21_X1  g540(.A(new_n565), .B1(new_n739), .B2(new_n377), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n728), .B(KEYINPUT51), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n377), .A2(new_n565), .A3(new_n606), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT52), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n735), .B2(new_n744), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n742), .B2(new_n748), .ZN(G1337gat));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(G99gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n736), .A2(new_n686), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n739), .A2(new_n690), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n750), .ZN(G1338gat));
  AOI21_X1  g552(.A(new_n673), .B1(new_n482), .B2(new_n637), .ZN(new_n754));
  INV_X1    g553(.A(new_n674), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n354), .B(new_n738), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(G106gat), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n607), .A2(new_n353), .A3(G106gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT53), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n730), .B2(new_n734), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(G106gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n756), .B2(KEYINPUT111), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n675), .A2(new_n767), .A3(new_n354), .A4(new_n738), .ZN(new_n768));
  AOI211_X1 g567(.A(KEYINPUT112), .B(new_n764), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(G106gat), .A3(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(new_n764), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n761), .B1(new_n769), .B2(new_n774), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n595), .A2(new_n597), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n776), .B2(new_n558), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n558), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n595), .A2(new_n779), .A3(new_n597), .A4(new_n559), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n602), .B1(new_n598), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(KEYINPUT55), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n604), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n783), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n557), .A2(new_n786), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n527), .A2(new_n528), .A3(new_n526), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n509), .B1(new_n520), .B2(new_n508), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n542), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n555), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n607), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n637), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n786), .A2(new_n790), .A3(new_n792), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n637), .A2(new_n555), .A3(new_n796), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n621), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n638), .A2(new_n667), .A3(new_n607), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n420), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(new_n376), .A3(new_n465), .ZN(new_n807));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n557), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n354), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n377), .A2(new_n420), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n686), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n811), .A2(new_n257), .A3(new_n667), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n808), .A2(new_n812), .ZN(G1340gat));
  NAND3_X1  g612(.A1(new_n807), .A2(new_n255), .A3(new_n606), .ZN(new_n814));
  OAI21_X1  g613(.A(G120gat), .B1(new_n811), .B2(new_n607), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT116), .Z(G1341gat));
  NAND3_X1  g616(.A1(new_n807), .A2(new_n250), .A3(new_n620), .ZN(new_n818));
  OAI21_X1  g617(.A(G127gat), .B1(new_n811), .B2(new_n621), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n663), .A2(new_n377), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n252), .A3(new_n465), .A4(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n811), .B2(new_n663), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G1343gat));
  NOR2_X1   g625(.A1(new_n690), .A2(new_n353), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT119), .Z(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n376), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n667), .A2(G141gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833));
  INV_X1    g632(.A(new_n805), .ZN(new_n834));
  XOR2_X1   g633(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n781), .B2(new_n783), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n785), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n798), .B1(new_n838), .B2(new_n557), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n637), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n604), .A3(new_n784), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n799), .B1(new_n667), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n803), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n834), .B1(new_n848), .B2(new_n621), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT57), .B1(new_n849), .B2(new_n353), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n472), .A2(new_n810), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n804), .A2(new_n805), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n354), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G141gat), .B1(new_n855), .B2(new_n667), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n832), .A2(new_n833), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n806), .A2(new_n376), .A3(new_n827), .A4(new_n831), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n859), .B2(new_n833), .ZN(G1344gat));
  NAND3_X1  g659(.A1(new_n830), .A2(new_n327), .A3(new_n606), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n852), .A2(KEYINPUT57), .A3(new_n354), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n803), .B1(new_n841), .B2(new_n845), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n805), .B1(new_n866), .B2(new_n620), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n353), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT121), .B(new_n805), .C1(new_n866), .C2(new_n620), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n871), .B2(KEYINPUT122), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(KEYINPUT57), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n606), .B(new_n851), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n855), .A2(new_n607), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n327), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n861), .B1(new_n876), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n830), .A2(new_n319), .A3(new_n620), .ZN(new_n880));
  OAI21_X1  g679(.A(G155gat), .B1(new_n855), .B2(new_n621), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1346gat));
  NAND3_X1  g681(.A1(new_n829), .A2(new_n320), .A3(new_n821), .ZN(new_n883));
  OAI21_X1  g682(.A(G162gat), .B1(new_n855), .B2(new_n663), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n376), .A2(new_n421), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n720), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n809), .A2(new_n557), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT123), .B1(new_n888), .B2(G169gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n421), .B1(new_n804), .B2(new_n805), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n377), .A3(new_n465), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n557), .A2(new_n237), .A3(new_n239), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n889), .A2(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT124), .ZN(G1348gat));
  NAND2_X1  g694(.A1(new_n809), .A2(new_n887), .ZN(new_n896));
  OAI21_X1  g695(.A(G176gat), .B1(new_n896), .B2(new_n607), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n606), .A2(new_n205), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n892), .B2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n896), .B2(new_n621), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n620), .A2(new_n212), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n900), .B(new_n901), .C1(new_n892), .C2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n896), .B2(new_n663), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n637), .A2(new_n213), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n892), .B2(new_n908), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n690), .A2(new_n376), .A3(new_n353), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n557), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n472), .A2(new_n886), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n863), .B(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n869), .A2(new_n870), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n853), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(new_n873), .ZN(new_n918));
  INV_X1    g717(.A(new_n874), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n557), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(new_n914), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n872), .B2(new_n874), .ZN(new_n924));
  OAI21_X1  g723(.A(G204gat), .B1(new_n924), .B2(new_n607), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n911), .A2(G204gat), .A3(new_n607), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n308), .A3(new_n620), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n620), .B(new_n923), .C1(new_n872), .C2(new_n874), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n912), .B2(new_n637), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n637), .A2(G218gat), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n920), .B2(KEYINPUT126), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n924), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n937), .B2(new_n939), .ZN(G1355gat));
endmodule


