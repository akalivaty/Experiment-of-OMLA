

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n691), .A2(n586), .ZN(n661) );
  NOR2_X1 U552 ( .A1(G2104), .A2(n522), .ZN(n866) );
  AND2_X1 U553 ( .A1(n527), .A2(n526), .ZN(G164) );
  AND2_X1 U554 ( .A1(n862), .A2(G102), .ZN(n516) );
  OR2_X1 U555 ( .A1(n690), .A2(n689), .ZN(n517) );
  AND2_X1 U556 ( .A1(n1003), .A2(n738), .ZN(n518) );
  XNOR2_X1 U557 ( .A(n590), .B(KEYINPUT100), .ZN(n591) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n685), .ZN(n589) );
  AND2_X1 U559 ( .A1(n655), .A2(n660), .ZN(n656) );
  NOR2_X1 U560 ( .A1(n725), .A2(n518), .ZN(n726) );
  NOR2_X1 U561 ( .A1(G651), .A2(n577), .ZN(n771) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U563 ( .A(KEYINPUT17), .B(n519), .Z(n861) );
  NAND2_X1 U564 ( .A1(G138), .A2(n861), .ZN(n520) );
  XNOR2_X1 U565 ( .A(KEYINPUT89), .B(n520), .ZN(n521) );
  INV_X1 U566 ( .A(G2105), .ZN(n522) );
  AND2_X1 U567 ( .A1(n522), .A2(G2104), .ZN(n862) );
  NOR2_X1 U568 ( .A1(n521), .A2(n516), .ZN(n527) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n865) );
  NAND2_X1 U570 ( .A1(G114), .A2(n865), .ZN(n524) );
  NAND2_X1 U571 ( .A1(G126), .A2(n866), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT88), .B(n525), .Z(n526) );
  NAND2_X1 U574 ( .A1(n865), .A2(G113), .ZN(n530) );
  NAND2_X1 U575 ( .A1(G101), .A2(n862), .ZN(n528) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U578 ( .A1(G125), .A2(n866), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G137), .A2(n861), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n775) );
  NAND2_X1 U583 ( .A1(n775), .A2(G86), .ZN(n535) );
  XOR2_X1 U584 ( .A(KEYINPUT77), .B(n535), .Z(n538) );
  INV_X1 U585 ( .A(G651), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G543), .A2(n540), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n536), .Z(n770) );
  NAND2_X1 U588 ( .A1(n770), .A2(G61), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U590 ( .A(KEYINPUT78), .B(n539), .ZN(n543) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NOR2_X1 U592 ( .A1(n577), .A2(n540), .ZN(n774) );
  NAND2_X1 U593 ( .A1(n774), .A2(G73), .ZN(n541) );
  XOR2_X1 U594 ( .A(KEYINPUT2), .B(n541), .Z(n542) );
  NOR2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n771), .A2(G48), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(G305) );
  NAND2_X1 U598 ( .A1(G63), .A2(n770), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G51), .A2(n771), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U601 ( .A(KEYINPUT6), .B(n548), .ZN(n555) );
  NAND2_X1 U602 ( .A1(n775), .A2(G89), .ZN(n549) );
  XNOR2_X1 U603 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G76), .A2(n774), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT5), .B(n552), .ZN(n553) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n553), .ZN(n554) );
  NOR2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(n556), .Z(G168) );
  NAND2_X1 U610 ( .A1(G64), .A2(n770), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G52), .A2(n771), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U613 ( .A1(G77), .A2(n774), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G90), .A2(n775), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U617 ( .A1(n563), .A2(n562), .ZN(G171) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(n564) );
  XNOR2_X1 U619 ( .A(KEYINPUT70), .B(n564), .ZN(G286) );
  NAND2_X1 U620 ( .A1(G50), .A2(n771), .ZN(n571) );
  NAND2_X1 U621 ( .A1(G62), .A2(n770), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G88), .A2(n775), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U624 ( .A1(G75), .A2(n774), .ZN(n567) );
  XNOR2_X1 U625 ( .A(KEYINPUT79), .B(n567), .ZN(n568) );
  NOR2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT80), .ZN(G303) );
  NAND2_X1 U629 ( .A1(G49), .A2(n771), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U632 ( .A1(n770), .A2(n575), .ZN(n576) );
  XNOR2_X1 U633 ( .A(n576), .B(KEYINPUT76), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G72), .A2(n774), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G85), .A2(n775), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U639 ( .A1(G60), .A2(n770), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G47), .A2(n771), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U642 ( .A1(n585), .A2(n584), .ZN(G290) );
  NOR2_X1 U643 ( .A1(G164), .A2(G1384), .ZN(n691) );
  NAND2_X1 U644 ( .A1(G160), .A2(G40), .ZN(n692) );
  INV_X1 U645 ( .A(n692), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G8), .A2(n661), .ZN(n685) );
  NOR2_X1 U647 ( .A1(G1981), .A2(G305), .ZN(n587) );
  XOR2_X1 U648 ( .A(n587), .B(KEYINPUT24), .Z(n588) );
  NOR2_X1 U649 ( .A1(n685), .A2(n588), .ZN(n690) );
  INV_X1 U650 ( .A(n589), .ZN(n655) );
  NOR2_X1 U651 ( .A1(G2084), .A2(n661), .ZN(n657) );
  NOR2_X1 U652 ( .A1(n657), .A2(n589), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(G8), .ZN(n592) );
  XNOR2_X1 U654 ( .A(KEYINPUT30), .B(n592), .ZN(n593) );
  NOR2_X1 U655 ( .A1(n593), .A2(G168), .ZN(n598) );
  XOR2_X1 U656 ( .A(KEYINPUT25), .B(G2078), .Z(n934) );
  NOR2_X1 U657 ( .A1(n934), .A2(n661), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT97), .ZN(n596) );
  INV_X1 U659 ( .A(G1961), .ZN(n995) );
  NAND2_X1 U660 ( .A1(n995), .A2(n661), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n601) );
  NOR2_X1 U662 ( .A1(G171), .A2(n601), .ZN(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U664 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n600), .B(n599), .ZN(n654) );
  NAND2_X1 U666 ( .A1(n601), .A2(G171), .ZN(n652) );
  INV_X1 U667 ( .A(n661), .ZN(n629) );
  NAND2_X1 U668 ( .A1(n629), .A2(G2072), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(KEYINPUT27), .ZN(n604) );
  AND2_X1 U670 ( .A1(G1956), .A2(n661), .ZN(n603) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n612) );
  NAND2_X1 U672 ( .A1(G65), .A2(n770), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G78), .A2(n774), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U675 ( .A1(G91), .A2(n775), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G53), .A2(n771), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n784) );
  NOR2_X1 U679 ( .A1(n612), .A2(n784), .ZN(n611) );
  XOR2_X1 U680 ( .A(n611), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U681 ( .A1(n612), .A2(n784), .ZN(n647) );
  NAND2_X1 U682 ( .A1(n770), .A2(G56), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT14), .B(n613), .Z(n621) );
  NAND2_X1 U684 ( .A1(n775), .A2(G81), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT12), .B(n614), .Z(n617) );
  NAND2_X1 U686 ( .A1(n774), .A2(G68), .ZN(n615) );
  XOR2_X1 U687 ( .A(n615), .B(KEYINPUT66), .Z(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT67), .B(n618), .Z(n619) );
  XNOR2_X1 U690 ( .A(n619), .B(KEYINPUT13), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n771), .A2(G43), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n982) );
  XOR2_X1 U694 ( .A(G1996), .B(KEYINPUT98), .Z(n935) );
  NOR2_X1 U695 ( .A1(n661), .A2(n935), .ZN(n625) );
  XOR2_X1 U696 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n661), .A2(G1341), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT99), .ZN(n641) );
  NAND2_X1 U701 ( .A1(G1348), .A2(n661), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G2067), .A2(n629), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n643) );
  NAND2_X1 U704 ( .A1(n771), .A2(G54), .ZN(n638) );
  NAND2_X1 U705 ( .A1(G66), .A2(n770), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G92), .A2(n775), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n774), .A2(G79), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT68), .B(n634), .Z(n635) );
  NOR2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT15), .B(n639), .Z(n997) );
  NAND2_X1 U713 ( .A1(n643), .A2(n997), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n982), .A2(n642), .ZN(n645) );
  NOR2_X1 U716 ( .A1(n643), .A2(n997), .ZN(n644) );
  NOR2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U720 ( .A(KEYINPUT29), .B(n650), .Z(n651) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n656), .B(KEYINPUT102), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n657), .A2(G8), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n670) );
  NAND2_X1 U726 ( .A1(G286), .A2(n660), .ZN(n666) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n685), .ZN(n663) );
  NOR2_X1 U728 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n664), .A2(G303), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(G8), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT32), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n683) );
  NOR2_X1 U735 ( .A1(G1976), .A2(G288), .ZN(n676) );
  NOR2_X1 U736 ( .A1(G303), .A2(G1971), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n676), .A2(n671), .ZN(n984) );
  NAND2_X1 U738 ( .A1(n683), .A2(n984), .ZN(n673) );
  NAND2_X1 U739 ( .A1(G288), .A2(G1976), .ZN(n672) );
  XOR2_X1 U740 ( .A(KEYINPUT103), .B(n672), .Z(n983) );
  NAND2_X1 U741 ( .A1(n673), .A2(n983), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n685), .A2(n674), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n675), .A2(KEYINPUT33), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n676), .A2(KEYINPUT33), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n677), .A2(n685), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U747 ( .A(G1981), .B(G305), .Z(n991) );
  NAND2_X1 U748 ( .A1(n680), .A2(n991), .ZN(n688) );
  NOR2_X1 U749 ( .A1(G303), .A2(G2090), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(KEYINPUT104), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n682), .A2(G8), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n693), .B(KEYINPUT90), .ZN(n738) );
  INV_X1 U757 ( .A(n738), .ZN(n714) );
  NAND2_X1 U758 ( .A1(n862), .A2(G105), .ZN(n695) );
  XNOR2_X1 U759 ( .A(KEYINPUT38), .B(KEYINPUT94), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n695), .B(n694), .ZN(n702) );
  NAND2_X1 U761 ( .A1(G117), .A2(n865), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G141), .A2(n861), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U764 ( .A1(G129), .A2(n866), .ZN(n698) );
  XNOR2_X1 U765 ( .A(KEYINPUT93), .B(n698), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n859) );
  NAND2_X1 U768 ( .A1(G1996), .A2(n859), .ZN(n712) );
  NAND2_X1 U769 ( .A1(G131), .A2(n861), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G95), .A2(n862), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT92), .B(n705), .ZN(n708) );
  NAND2_X1 U773 ( .A1(G107), .A2(n865), .ZN(n706) );
  XNOR2_X1 U774 ( .A(KEYINPUT91), .B(n706), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U776 ( .A1(n866), .A2(G119), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n879) );
  NAND2_X1 U778 ( .A1(G1991), .A2(n879), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(KEYINPUT95), .B(n713), .ZN(n959) );
  NOR2_X1 U781 ( .A1(n714), .A2(n959), .ZN(n730) );
  XOR2_X1 U782 ( .A(KEYINPUT96), .B(n730), .Z(n724) );
  XNOR2_X1 U783 ( .A(G2067), .B(KEYINPUT37), .ZN(n735) );
  NAND2_X1 U784 ( .A1(G116), .A2(n865), .ZN(n716) );
  NAND2_X1 U785 ( .A1(G128), .A2(n866), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U787 ( .A(n717), .B(KEYINPUT35), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G140), .A2(n861), .ZN(n719) );
  NAND2_X1 U789 ( .A1(G104), .A2(n862), .ZN(n718) );
  NAND2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U791 ( .A(KEYINPUT34), .B(n720), .Z(n721) );
  NAND2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U793 ( .A(n723), .B(KEYINPUT36), .Z(n872) );
  NOR2_X1 U794 ( .A1(n735), .A2(n872), .ZN(n963) );
  NAND2_X1 U795 ( .A1(n963), .A2(n738), .ZN(n733) );
  NAND2_X1 U796 ( .A1(n724), .A2(n733), .ZN(n725) );
  XNOR2_X1 U797 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U798 ( .A1(n517), .A2(n726), .ZN(n741) );
  NOR2_X1 U799 ( .A1(G1996), .A2(n859), .ZN(n956) );
  NOR2_X1 U800 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U801 ( .A1(G1991), .A2(n879), .ZN(n962) );
  NOR2_X1 U802 ( .A1(n727), .A2(n962), .ZN(n728) );
  XOR2_X1 U803 ( .A(KEYINPUT105), .B(n728), .Z(n729) );
  NOR2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n956), .A2(n731), .ZN(n732) );
  XNOR2_X1 U806 ( .A(KEYINPUT39), .B(n732), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n734), .A2(n733), .ZN(n737) );
  AND2_X1 U808 ( .A1(n735), .A2(n872), .ZN(n736) );
  XOR2_X1 U809 ( .A(KEYINPUT106), .B(n736), .Z(n973) );
  NAND2_X1 U810 ( .A1(n737), .A2(n973), .ZN(n739) );
  NAND2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U813 ( .A(n742), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U814 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U815 ( .A(G132), .ZN(G219) );
  INV_X1 U816 ( .A(G120), .ZN(G236) );
  INV_X1 U817 ( .A(G69), .ZN(G235) );
  INV_X1 U818 ( .A(G57), .ZN(G237) );
  INV_X1 U819 ( .A(n784), .ZN(G299) );
  NAND2_X1 U820 ( .A1(G7), .A2(G661), .ZN(n743) );
  XNOR2_X1 U821 ( .A(n743), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U822 ( .A(G223), .ZN(n813) );
  NAND2_X1 U823 ( .A1(n813), .A2(G567), .ZN(n744) );
  XOR2_X1 U824 ( .A(KEYINPUT11), .B(n744), .Z(G234) );
  INV_X1 U825 ( .A(G860), .ZN(n750) );
  OR2_X1 U826 ( .A1(n982), .A2(n750), .ZN(G153) );
  INV_X1 U827 ( .A(G171), .ZN(G301) );
  NAND2_X1 U828 ( .A1(G868), .A2(G301), .ZN(n746) );
  INV_X1 U829 ( .A(G868), .ZN(n793) );
  NAND2_X1 U830 ( .A1(n997), .A2(n793), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(G284) );
  XNOR2_X1 U832 ( .A(KEYINPUT71), .B(G868), .ZN(n747) );
  NOR2_X1 U833 ( .A1(G286), .A2(n747), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G868), .A2(G299), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n749), .A2(n748), .ZN(G297) );
  NAND2_X1 U836 ( .A1(n750), .A2(G559), .ZN(n751) );
  INV_X1 U837 ( .A(n997), .ZN(n885) );
  NAND2_X1 U838 ( .A1(n751), .A2(n885), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT16), .ZN(n753) );
  XNOR2_X1 U840 ( .A(KEYINPUT72), .B(n753), .ZN(G148) );
  NOR2_X1 U841 ( .A1(n997), .A2(n793), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n754), .B(KEYINPUT73), .ZN(n755) );
  NOR2_X1 U843 ( .A1(G559), .A2(n755), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT74), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n982), .A2(G868), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(G282) );
  NAND2_X1 U847 ( .A1(G111), .A2(n865), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G99), .A2(n862), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n766) );
  NAND2_X1 U850 ( .A1(n866), .A2(G123), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT18), .ZN(n763) );
  NAND2_X1 U852 ( .A1(G135), .A2(n861), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U854 ( .A(KEYINPUT75), .B(n764), .Z(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n961) );
  XNOR2_X1 U856 ( .A(n961), .B(G2096), .ZN(n768) );
  INV_X1 U857 ( .A(G2100), .ZN(n767) );
  NAND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(G156) );
  NAND2_X1 U859 ( .A1(n885), .A2(G559), .ZN(n791) );
  XNOR2_X1 U860 ( .A(n982), .B(n791), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n769), .A2(G860), .ZN(n780) );
  NAND2_X1 U862 ( .A1(G67), .A2(n770), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G55), .A2(n771), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G80), .A2(n774), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G93), .A2(n775), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n794) );
  XNOR2_X1 U869 ( .A(n780), .B(n794), .ZN(G145) );
  XOR2_X1 U870 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n782) );
  XNOR2_X1 U871 ( .A(KEYINPUT83), .B(KEYINPUT81), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n794), .B(n783), .ZN(n786) );
  XNOR2_X1 U874 ( .A(G290), .B(n784), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U876 ( .A(n787), .B(G305), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n788), .B(G288), .ZN(n789) );
  XNOR2_X1 U878 ( .A(G303), .B(n789), .ZN(n790) );
  XNOR2_X1 U879 ( .A(n790), .B(n982), .ZN(n884) );
  XOR2_X1 U880 ( .A(n884), .B(n791), .Z(n792) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n796) );
  NOR2_X1 U882 ( .A1(G868), .A2(n794), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U884 ( .A(KEYINPUT84), .B(n797), .Z(G295) );
  NAND2_X1 U885 ( .A1(G2084), .A2(G2078), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT20), .B(n798), .Z(n799) );
  NAND2_X1 U887 ( .A1(G2090), .A2(n799), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT21), .B(n800), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n801), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U890 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U891 ( .A(KEYINPUT65), .B(G82), .ZN(G220) );
  NOR2_X1 U892 ( .A1(G235), .A2(G236), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n802), .B(KEYINPUT85), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G237), .A2(n803), .ZN(n804) );
  XNOR2_X1 U895 ( .A(KEYINPUT86), .B(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n805), .A2(G108), .ZN(n817) );
  NAND2_X1 U897 ( .A1(n817), .A2(G567), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G219), .A2(G220), .ZN(n806) );
  XOR2_X1 U899 ( .A(KEYINPUT22), .B(n806), .Z(n807) );
  NOR2_X1 U900 ( .A1(G218), .A2(n807), .ZN(n808) );
  NAND2_X1 U901 ( .A1(G96), .A2(n808), .ZN(n818) );
  NAND2_X1 U902 ( .A1(n818), .A2(G2106), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G483), .A2(G661), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n819), .A2(n811), .ZN(n812) );
  XOR2_X1 U906 ( .A(KEYINPUT87), .B(n812), .Z(n816) );
  NAND2_X1 U907 ( .A1(n816), .A2(G36), .ZN(G176) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U910 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(G188) );
  XOR2_X1 U913 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  NOR2_X1 U916 ( .A1(n818), .A2(n817), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  INV_X1 U918 ( .A(n819), .ZN(G319) );
  XNOR2_X1 U919 ( .A(G1991), .B(KEYINPUT41), .ZN(n829) );
  XOR2_X1 U920 ( .A(G1976), .B(G1971), .Z(n821) );
  XNOR2_X1 U921 ( .A(G1996), .B(G1961), .ZN(n820) );
  XNOR2_X1 U922 ( .A(n821), .B(n820), .ZN(n825) );
  XOR2_X1 U923 ( .A(G1981), .B(G1956), .Z(n823) );
  XNOR2_X1 U924 ( .A(G1986), .B(G1966), .ZN(n822) );
  XNOR2_X1 U925 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U926 ( .A(n825), .B(n824), .Z(n827) );
  XNOR2_X1 U927 ( .A(KEYINPUT114), .B(G2474), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(G229) );
  XOR2_X1 U930 ( .A(G2096), .B(G2090), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2084), .B(G2072), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U933 ( .A(KEYINPUT109), .B(KEYINPUT113), .Z(n833) );
  XNOR2_X1 U934 ( .A(G2100), .B(KEYINPUT110), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n842) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2678), .B(KEYINPUT42), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n838), .B(KEYINPUT111), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2078), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(G227) );
  NAND2_X1 U944 ( .A1(G124), .A2(n866), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n843), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G136), .A2(n861), .ZN(n844) );
  XOR2_X1 U947 ( .A(KEYINPUT115), .B(n844), .Z(n845) );
  NAND2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U949 ( .A1(G112), .A2(n865), .ZN(n848) );
  NAND2_X1 U950 ( .A1(G100), .A2(n862), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U952 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U953 ( .A1(G142), .A2(n861), .ZN(n852) );
  NAND2_X1 U954 ( .A1(G106), .A2(n862), .ZN(n851) );
  NAND2_X1 U955 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT45), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G118), .A2(n865), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G130), .A2(n866), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT116), .B(n856), .Z(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n877) );
  NAND2_X1 U963 ( .A1(G139), .A2(n861), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G103), .A2(n862), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G115), .A2(n865), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G127), .A2(n866), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n966) );
  XOR2_X1 U971 ( .A(n961), .B(G162), .Z(n874) );
  XOR2_X1 U972 ( .A(G164), .B(n872), .Z(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(n966), .B(n875), .Z(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n882) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U978 ( .A(G160), .B(n880), .Z(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U980 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U981 ( .A(n884), .B(KEYINPUT117), .ZN(n887) );
  XNOR2_X1 U982 ( .A(G171), .B(n885), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(G286), .ZN(n889) );
  NOR2_X1 U985 ( .A1(G37), .A2(n889), .ZN(G397) );
  XNOR2_X1 U986 ( .A(G2443), .B(G2427), .ZN(n899) );
  XOR2_X1 U987 ( .A(G2430), .B(KEYINPUT108), .Z(n891) );
  XNOR2_X1 U988 ( .A(G2454), .B(G2435), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U990 ( .A(G2438), .B(KEYINPUT107), .Z(n893) );
  XNOR2_X1 U991 ( .A(G1348), .B(G1341), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2451), .B(G2446), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n900), .A2(G14), .ZN(n906) );
  NAND2_X1 U998 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(n906), .ZN(G401) );
  INV_X1 U1006 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1007 ( .A(G5), .B(n995), .ZN(n920) );
  XNOR2_X1 U1008 ( .A(G1966), .B(G21), .ZN(n918) );
  XNOR2_X1 U1009 ( .A(G1956), .B(G20), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n907), .B(G4), .ZN(n908) );
  XNOR2_X1 U1012 ( .A(n908), .B(G1348), .ZN(n909) );
  NOR2_X1 U1013 ( .A1(n910), .A2(n909), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G19), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(G1981), .B(G6), .ZN(n911) );
  NOR2_X1 U1016 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(n915), .B(KEYINPUT60), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(KEYINPUT126), .B(n916), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(G1986), .B(G24), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(G22), .B(G1971), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G1976), .B(KEYINPUT127), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(n923), .B(G23), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n926), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1030 ( .A(KEYINPUT61), .B(n929), .Z(n930) );
  NOR2_X1 U1031 ( .A1(G16), .A2(n930), .ZN(n954) );
  XNOR2_X1 U1032 ( .A(G1991), .B(G25), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n941) );
  XOR2_X1 U1035 ( .A(G2067), .B(G26), .Z(n933) );
  NAND2_X1 U1036 ( .A1(n933), .A2(G28), .ZN(n939) );
  XOR2_X1 U1037 ( .A(n934), .B(G27), .Z(n937) );
  XNOR2_X1 U1038 ( .A(n935), .B(G32), .ZN(n936) );
  NAND2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(KEYINPUT53), .ZN(n945) );
  XOR2_X1 U1043 ( .A(G2084), .B(G34), .Z(n943) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(n943), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(KEYINPUT55), .B(n948), .ZN(n950) );
  INV_X1 U1049 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(n951), .A2(G11), .ZN(n952) );
  XOR2_X1 U1052 ( .A(KEYINPUT119), .B(n952), .Z(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n981) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1056 ( .A(KEYINPUT51), .B(n957), .Z(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n975) );
  XOR2_X1 U1058 ( .A(G2084), .B(G160), .Z(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n971) );
  XOR2_X1 U1062 ( .A(G2072), .B(n966), .Z(n968) );
  XOR2_X1 U1063 ( .A(G164), .B(G2078), .Z(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1065 ( .A(KEYINPUT50), .B(n969), .Z(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n976), .ZN(n978) );
  INV_X1 U1070 ( .A(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n979), .A2(G29), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n1013) );
  XOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .Z(n1010) );
  XOR2_X1 U1075 ( .A(n982), .B(G1341), .Z(n990) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n987) );
  INV_X1 U1077 ( .A(G1971), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(G166), .A2(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n988), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1007) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT57), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT120), .B(n994), .ZN(n1005) );
  XNOR2_X1 U1086 ( .A(n995), .B(G171), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT121), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G299), .B(G1956), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n997), .B(G1348), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT123), .B(n1008), .Z(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1011), .B(KEYINPUT124), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1014), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

