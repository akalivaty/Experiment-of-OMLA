//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  OR2_X1    g000(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT64), .A2(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G146), .A3(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n189), .A2(new_n194), .A3(new_n199), .A4(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(G143), .B1(new_n191), .B2(new_n193), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n197), .B2(new_n198), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n187), .A2(new_n188), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n194), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n200), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G137), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n208), .A2(G137), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n208), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n209), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n209), .A3(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n218), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n194), .A2(new_n199), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n201), .B2(new_n202), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT2), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT2), .A3(G113), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n234), .A2(new_n236), .B1(new_n232), .B2(new_n233), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(G116), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n240), .A2(KEYINPUT69), .A3(new_n241), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n240), .B2(new_n241), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n237), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n221), .A3(new_n230), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n260), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n258), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n256), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT65), .B(G146), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(G143), .B1(new_n187), .B2(new_n188), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n271), .A2(new_n204), .B1(new_n202), .B2(new_n201), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n219), .B1(new_n272), .B2(new_n200), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n230), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n225), .A2(new_n227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n192), .A2(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n196), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT64), .A2(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT64), .A2(G143), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n190), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n276), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n194), .A2(new_n199), .A3(new_n225), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT66), .A3(new_n224), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n273), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT71), .B1(new_n287), .B2(new_n249), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT66), .B1(new_n285), .B2(new_n224), .ZN(new_n289));
  AND4_X1   g103(.A1(KEYINPUT66), .A2(new_n224), .A3(new_n226), .A4(new_n229), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n221), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n247), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n293), .A3(new_n250), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT28), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n258), .A2(new_n267), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(KEYINPUT72), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n221), .A2(KEYINPUT30), .A3(new_n230), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n247), .B(new_n298), .C1(new_n287), .C2(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n250), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n300), .B2(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT72), .B1(new_n295), .B2(new_n296), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n269), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G472), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n266), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n250), .A3(new_n266), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT31), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n299), .A2(new_n311), .A3(new_n250), .A4(new_n266), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(KEYINPUT32), .B(new_n306), .C1(new_n308), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n258), .B1(new_n294), .B2(KEYINPUT28), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n310), .B(new_n312), .C1(new_n317), .C2(new_n266), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n306), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n306), .B1(new_n308), .B2(new_n313), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n305), .A2(new_n316), .A3(new_n319), .A4(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT9), .B(G234), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT79), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G902), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G221), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT80), .Z(new_n330));
  INV_X1    g144(.A(G469), .ZN(new_n331));
  INV_X1    g145(.A(new_n224), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G104), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(KEYINPUT3), .A3(G107), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n336), .A2(KEYINPUT82), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n337), .B1(new_n342), .B2(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(KEYINPUT82), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(G104), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G107), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT83), .A4(G107), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n194), .A2(new_n199), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n204), .B1(new_n282), .B2(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n200), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n342), .B1(G104), .B2(new_n338), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n207), .B1(new_n352), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n335), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n333), .A2(new_n334), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n343), .A2(new_n350), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G101), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n351), .B1(new_n343), .B2(new_n350), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n285), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n352), .A2(new_n207), .A3(KEYINPUT10), .A4(new_n357), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n368), .A2(new_n332), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  OAI221_X1 g187(.A(new_n335), .B1(new_n333), .B2(new_n334), .C1(new_n358), .C2(new_n359), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT81), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n262), .A2(G227), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND4_X1  g192(.A1(new_n362), .A2(new_n373), .A3(new_n374), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n366), .A2(new_n367), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n365), .A2(new_n285), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n369), .B(new_n372), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n224), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n378), .B1(new_n383), .B2(new_n373), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g200(.A(KEYINPUT85), .B(new_n378), .C1(new_n383), .C2(new_n373), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n331), .B(new_n327), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n362), .A2(new_n373), .A3(new_n374), .ZN(new_n389));
  INV_X1    g203(.A(new_n378), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n383), .A2(new_n378), .A3(new_n373), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(G469), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n331), .A2(new_n327), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n330), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n247), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n400));
  INV_X1    g214(.A(new_n243), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT5), .B1(new_n244), .B2(new_n245), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n233), .B1(new_n403), .B2(new_n239), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n405), .B2(KEYINPUT86), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n406), .A2(new_n352), .A3(new_n357), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n400), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n409), .A3(new_n411), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G125), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n272), .A2(new_n416), .A3(new_n200), .ZN(new_n417));
  OAI21_X1  g231(.A(G125), .B1(new_n283), .B2(new_n284), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G224), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G953), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n423), .A3(new_n412), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT7), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(new_n420), .B2(G953), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n417), .A2(new_n418), .A3(new_n429), .A4(new_n427), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n404), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n352), .B(new_n357), .C1(new_n401), .C2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n411), .B(KEYINPUT8), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n406), .A2(new_n408), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n352), .A2(new_n357), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n414), .A2(new_n433), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n441), .A2(new_n327), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n425), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n425), .A2(new_n444), .A3(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n399), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n397), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n416), .A2(G140), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT16), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n450), .A3(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G146), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n190), .A2(KEYINPUT75), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(G146), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n453), .A2(new_n455), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n261), .A2(new_n262), .A3(G214), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n197), .A3(new_n198), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n261), .A2(new_n262), .A3(G143), .A4(G214), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n217), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n458), .A2(new_n461), .B1(new_n465), .B2(KEYINPUT17), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n217), .A3(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(KEYINPUT17), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT89), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n336), .ZN(new_n474));
  XNOR2_X1  g288(.A(G125), .B(G140), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n270), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n190), .B2(new_n475), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT18), .A2(G131), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n464), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n465), .A2(KEYINPUT18), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n471), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n474), .B1(new_n471), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G475), .B1(new_n486), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n489));
  INV_X1    g303(.A(new_n469), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n465), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n468), .A2(KEYINPUT88), .A3(new_n469), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n453), .A2(G146), .A3(new_n455), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n475), .B(KEYINPUT19), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n270), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n493), .A2(new_n497), .B1(new_n481), .B2(new_n480), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n483), .B1(new_n498), .B2(new_n474), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(KEYINPUT90), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n499), .A2(new_n505), .A3(new_n500), .A4(new_n501), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n488), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(G952), .A3(new_n262), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT99), .Z(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(G902), .A3(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT21), .B(G898), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n517));
  INV_X1    g331(.A(G122), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G116), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n238), .A2(G122), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n238), .A2(G122), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(G116), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT91), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n338), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(G107), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n197), .A2(G128), .A3(new_n198), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT13), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n196), .A2(G128), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI221_X1 g348(.A(G134), .B1(new_n529), .B2(new_n530), .C1(new_n531), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(new_n208), .A3(new_n533), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(KEYINPUT93), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(KEYINPUT93), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n528), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n540));
  AOI21_X1  g354(.A(G107), .B1(new_n521), .B2(new_n524), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n518), .B2(G116), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT94), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n522), .A2(new_n544), .A3(KEYINPUT14), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n518), .A2(KEYINPUT14), .A3(G116), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n523), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(G107), .B2(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n280), .A2(new_n281), .A3(new_n204), .ZN(new_n549));
  OAI21_X1  g363(.A(G134), .B1(new_n549), .B2(new_n532), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n536), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n540), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(G107), .ZN(new_n553));
  AND4_X1   g367(.A1(new_n540), .A2(new_n551), .A3(new_n526), .A4(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n539), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G217), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n325), .A2(new_n556), .A3(G953), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n539), .B(new_n557), .C1(new_n552), .C2(new_n554), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT96), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n562), .A3(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n327), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G478), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n564), .A2(new_n565), .A3(new_n567), .A4(G478), .ZN(new_n570));
  AND4_X1   g384(.A1(KEYINPUT97), .A2(new_n561), .A3(new_n327), .A4(new_n563), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT98), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n568), .B2(new_n566), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n570), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n516), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n239), .B2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n239), .A2(G128), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(G119), .B(G128), .ZN(new_n584));
  INV_X1    g398(.A(G110), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT24), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT24), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G110), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n583), .A2(G110), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n458), .A2(new_n461), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n458), .A2(new_n590), .A3(new_n593), .A4(new_n461), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n494), .A2(new_n476), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n580), .A2(new_n582), .A3(new_n585), .A4(new_n581), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT77), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n204), .A2(G119), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n581), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT24), .B(G110), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n597), .A2(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n596), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n595), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT78), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT22), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n215), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(KEYINPUT25), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n556), .B1(G234), .B2(new_n327), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n613), .A2(new_n615), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT25), .B1(new_n621), .B2(G902), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT78), .B1(new_n595), .B2(new_n605), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n607), .B(new_n604), .C1(new_n592), .C2(new_n594), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n614), .B1(new_n625), .B2(new_n612), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n618), .A2(G902), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n620), .A2(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n323), .A2(new_n449), .A3(new_n578), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  AND3_X1   g444(.A1(new_n425), .A2(new_n444), .A3(new_n442), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n444), .B1(new_n425), .B2(new_n442), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n398), .B(new_n515), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n504), .A2(new_n506), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n487), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n561), .A2(new_n636), .A3(new_n563), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n559), .A2(KEYINPUT33), .A3(new_n560), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(G478), .A3(new_n327), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G478), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n564), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n633), .B2(new_n643), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n487), .A2(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n448), .A2(new_n645), .A3(new_n646), .A4(new_n515), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n327), .B1(new_n308), .B2(new_n313), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n318), .B(new_n327), .C1(new_n650), .C2(new_n651), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n628), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n388), .A2(new_n396), .ZN(new_n656));
  INV_X1    g470(.A(new_n330), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  AND2_X1   g476(.A1(new_n574), .A2(new_n577), .ZN(new_n663));
  INV_X1    g477(.A(new_n502), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n487), .B1(new_n664), .B2(new_n503), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n633), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n659), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  AND2_X1   g483(.A1(new_n653), .A2(new_n654), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n625), .B1(KEYINPUT36), .B2(new_n612), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n623), .B2(new_n624), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n627), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT25), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n626), .B2(new_n327), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n676), .B2(new_n619), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n679), .B(new_n674), .C1(new_n676), .C2(new_n619), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n449), .A2(new_n578), .A3(new_n670), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G110), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  NAND2_X1  g499(.A1(new_n446), .A2(new_n447), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n686), .A3(new_n398), .A4(new_n680), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n658), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n511), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n510), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n487), .B(new_n692), .C1(new_n664), .C2(new_n503), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n574), .A2(new_n577), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n695), .A3(new_n323), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n688), .A2(new_n695), .A3(new_n323), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XOR2_X1   g515(.A(new_n691), .B(KEYINPUT39), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n397), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT40), .Z(new_n704));
  INV_X1    g518(.A(new_n677), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n398), .A2(new_n663), .A3(new_n635), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n631), .A2(new_n632), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT38), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT38), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n316), .A2(new_n319), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT32), .B1(new_n318), .B2(new_n306), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n251), .A2(new_n267), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n309), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(G902), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(G472), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n704), .A2(new_n706), .A3(new_n713), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n197), .A2(new_n198), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G45));
  NOR2_X1   g538(.A1(new_n643), .A2(new_n691), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n688), .A2(new_n323), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  INV_X1    g541(.A(new_n628), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n716), .B1(G472), .B2(new_n304), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n715), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n327), .B1(new_n386), .B2(new_n387), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n329), .A3(new_n388), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n648), .A3(KEYINPUT106), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n256), .A2(new_n268), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n327), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n221), .A2(KEYINPUT30), .A3(new_n230), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n738), .B1(new_n291), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n257), .B1(new_n740), .B2(new_n247), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n259), .B1(new_n741), .B2(new_n266), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n307), .A2(new_n266), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n294), .B2(KEYINPUT28), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(new_n744), .B2(KEYINPUT72), .ZN(new_n745));
  INV_X1    g559(.A(new_n303), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n737), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n322), .B1(new_n747), .B2(new_n651), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n733), .B(new_n628), .C1(new_n748), .C2(new_n714), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n644), .A2(new_n647), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n735), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n734), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT41), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G113), .ZN(G15));
  NAND2_X1  g568(.A1(new_n663), .A2(new_n666), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n238), .ZN(G18));
  NAND3_X1  g571(.A1(new_n732), .A2(new_n329), .A3(new_n388), .ZN(new_n758));
  INV_X1    g572(.A(new_n448), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n323), .A3(new_n578), .A4(new_n681), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  AND4_X1   g576(.A1(new_n448), .A2(new_n574), .A3(new_n577), .A4(new_n635), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n649), .A2(G472), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n266), .B1(new_n256), .B2(new_n307), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n306), .B1(new_n765), .B2(new_n313), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n764), .A2(new_n628), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n758), .A2(new_n514), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  AND3_X1   g584(.A1(new_n764), .A2(new_n677), .A3(new_n766), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n760), .A2(new_n725), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n392), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n383), .A2(KEYINPUT107), .A3(new_n378), .A4(new_n373), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(G469), .A3(new_n391), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n388), .A2(new_n395), .A3(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n631), .A2(new_n632), .A3(new_n399), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n779), .A2(new_n329), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n323), .A2(new_n781), .A3(new_n628), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n725), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n774), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  INV_X1    g600(.A(new_n314), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT108), .B1(new_n787), .B2(new_n716), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n322), .A2(new_n789), .A3(new_n314), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n305), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n628), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(KEYINPUT109), .A3(new_n628), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n781), .A2(KEYINPUT42), .A3(new_n725), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n786), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n791), .A2(KEYINPUT109), .A3(new_n628), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT109), .B1(new_n791), .B2(new_n628), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n786), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n785), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND2_X1  g618(.A1(new_n782), .A2(new_n695), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  INV_X1    g620(.A(new_n780), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n635), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n507), .A2(KEYINPUT111), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n642), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT43), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n642), .A2(new_n813), .A3(new_n507), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n670), .A3(new_n705), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n807), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n391), .B2(new_n392), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n331), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n776), .A2(KEYINPUT45), .A3(new_n391), .A4(new_n777), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n394), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n388), .B1(new_n822), .B2(KEYINPUT46), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n329), .B(new_n702), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n818), .B(new_n826), .C1(new_n817), .C2(new_n816), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT112), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  OAI21_X1  g643(.A(new_n329), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT47), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT47), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n323), .A2(new_n784), .A3(new_n628), .A4(new_n807), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n732), .A2(new_n388), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n657), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n831), .B2(new_n832), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n815), .ZN(new_n841));
  INV_X1    g655(.A(new_n510), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n767), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n807), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n836), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n758), .A2(new_n807), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n841), .A2(new_n842), .A3(new_n771), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n721), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n628), .A3(new_n842), .A4(new_n846), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n507), .A2(new_n641), .A3(new_n639), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n841), .A2(new_n842), .A3(new_n733), .A4(new_n767), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n399), .B1(new_n711), .B2(new_n712), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n855), .A3(KEYINPUT50), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n852), .B2(new_n854), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n851), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n845), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n796), .A2(new_n842), .A3(new_n841), .A4(new_n846), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n849), .A2(new_n643), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n853), .B2(new_n448), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n840), .B2(new_n844), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n807), .A4(new_n843), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n867), .A2(new_n868), .B1(new_n859), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n859), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n836), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT118), .B(new_n836), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n865), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n778), .A2(new_n395), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n877), .A2(new_n388), .B1(G221), .B2(new_n328), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n771), .A2(new_n725), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n678), .A2(new_n680), .A3(new_n694), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n573), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n575), .A2(KEYINPUT113), .A3(new_n570), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n397), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n748), .A2(new_n714), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n886), .A2(new_n780), .B1(new_n782), .B2(new_n695), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n629), .A2(new_n682), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n756), .ZN(new_n889));
  INV_X1    g703(.A(new_n633), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n635), .B1(new_n882), .B2(new_n883), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n659), .B(new_n890), .C1(new_n645), .C2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n892), .A2(new_n761), .A3(new_n769), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n887), .A2(new_n889), .A3(new_n893), .A4(new_n752), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT110), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n801), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n785), .ZN(new_n898));
  INV_X1    g712(.A(new_n772), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n697), .B2(new_n699), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n726), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g716(.A(KEYINPUT114), .B(new_n899), .C1(new_n697), .C2(new_n699), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n878), .A2(new_n705), .A3(new_n692), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n721), .A3(new_n763), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT52), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n905), .A2(new_n726), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT52), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n898), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n900), .A2(new_n908), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT52), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n900), .A2(KEYINPUT52), .A3(new_n908), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n898), .A2(KEYINPUT53), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  INV_X1    g734(.A(new_n894), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n803), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n916), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n909), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n911), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT115), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n898), .B2(new_n917), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n898), .B(KEYINPUT53), .C1(new_n907), .C2(new_n909), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n876), .A2(new_n920), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(G952), .B(new_n262), .C1(new_n933), .C2(KEYINPUT119), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n713), .A2(new_n721), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n628), .A2(new_n657), .A3(new_n398), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n938), .B(new_n811), .C1(KEYINPUT49), .C2(new_n837), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n937), .B(new_n939), .C1(KEYINPUT49), .C2(new_n837), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n936), .A3(new_n940), .ZN(G75));
  NAND3_X1  g755(.A1(new_n926), .A2(new_n929), .A3(new_n931), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(G210), .A3(G902), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n415), .A2(new_n424), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n422), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT55), .Z(new_n947));
  AND3_X1   g761(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n943), .B2(new_n944), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n262), .A2(G952), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(G51));
  OAI21_X1  g765(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n952));
  AOI211_X1 g766(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n898), .C2(new_n917), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT54), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n932), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n394), .B(KEYINPUT57), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n387), .B2(new_n386), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n820), .A2(new_n821), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n942), .A2(G902), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n950), .B1(new_n958), .B2(new_n963), .ZN(G54));
  INV_X1    g778(.A(new_n499), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n942), .A2(G902), .ZN(new_n966));
  NAND2_X1  g780(.A1(KEYINPUT58), .A2(G475), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n950), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n966), .A2(new_n965), .A3(new_n967), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G60));
  NAND2_X1  g786(.A1(new_n637), .A2(new_n638), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n640), .A2(new_n327), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n955), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n979), .A3(new_n969), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n920), .A2(new_n932), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n973), .B1(new_n981), .B2(new_n976), .ZN(new_n982));
  INV_X1    g796(.A(new_n977), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n954), .B2(new_n932), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT122), .B1(new_n984), .B2(new_n950), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n980), .A2(new_n982), .A3(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n942), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n626), .B(KEYINPUT123), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n942), .A2(new_n673), .A3(new_n671), .A4(new_n989), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n969), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n969), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  NAND3_X1  g812(.A1(new_n889), .A2(new_n893), .A3(new_n752), .ZN(new_n999));
  NAND2_X1  g813(.A1(G224), .A2(G953), .ZN(new_n1000));
  OAI22_X1  g814(.A1(new_n999), .A2(G953), .B1(new_n512), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(G898), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n945), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G69));
  AOI21_X1  g818(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n740), .B(new_n496), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n689), .B2(new_n262), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n902), .B2(new_n903), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n700), .A2(new_n772), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT114), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n900), .A2(new_n901), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(KEYINPUT124), .A3(new_n726), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1009), .A2(new_n1013), .A3(new_n827), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT125), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1009), .A2(new_n1013), .A3(new_n1016), .A4(new_n827), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n796), .A2(new_n763), .A3(new_n826), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n803), .A2(new_n1018), .A3(new_n805), .A4(new_n834), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AND4_X1   g834(.A1(KEYINPUT126), .A2(new_n1015), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1019), .B1(new_n1014), .B2(KEYINPUT125), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT126), .B1(new_n1022), .B2(new_n1017), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1007), .B1(new_n1024), .B2(new_n262), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1009), .A2(new_n1013), .A3(new_n722), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n703), .A2(new_n807), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n730), .B(new_n1029), .C1(new_n645), .C2(new_n891), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n827), .A2(new_n834), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1027), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1006), .B1(new_n1032), .B2(new_n262), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1005), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1033), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1005), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1021), .A2(new_n1023), .A3(G953), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1035), .B(new_n1036), .C1(new_n1037), .C2(new_n1007), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1034), .A2(new_n1038), .ZN(G72));
  XNOR2_X1  g853(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n300), .A2(new_n267), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n309), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n919), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(new_n969), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1023), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1022), .A2(KEYINPUT126), .A3(new_n1017), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n300), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1042), .B1(new_n1049), .B2(new_n999), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n300), .A2(new_n1042), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1044), .B1(new_n1032), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1046), .B1(new_n1050), .B2(new_n1052), .ZN(G57));
endmodule


