

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n522), .B(n521), .ZN(n645) );
  OR2_X1 U551 ( .A1(n697), .A2(n696), .ZN(n794) );
  BUF_X1 U552 ( .A(n690), .Z(n612) );
  INV_X2 U553 ( .A(G2105), .ZN(n540) );
  XNOR2_X1 U554 ( .A(n734), .B(n733), .ZN(n735) );
  AND2_X1 U555 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U556 ( .A1(n580), .A2(n579), .ZN(n702) );
  OR2_X1 U557 ( .A1(n728), .A2(G301), .ZN(n516) );
  OR2_X1 U558 ( .A1(n772), .A2(n787), .ZN(n517) );
  NOR2_X1 U559 ( .A1(n826), .A2(n825), .ZN(n518) );
  XOR2_X1 U560 ( .A(KEYINPUT94), .B(KEYINPUT32), .Z(n519) );
  XOR2_X1 U561 ( .A(n739), .B(n738), .Z(n520) );
  AND2_X1 U562 ( .A1(n724), .A2(G1996), .ZN(n698) );
  INV_X1 U563 ( .A(KEYINPUT90), .ZN(n704) );
  INV_X1 U564 ( .A(KEYINPUT91), .ZN(n733) );
  INV_X1 U565 ( .A(KEYINPUT31), .ZN(n737) );
  XNOR2_X1 U566 ( .A(n737), .B(KEYINPUT93), .ZN(n738) );
  NOR2_X1 U567 ( .A1(G1966), .A2(n741), .ZN(n754) );
  NAND2_X1 U568 ( .A1(n795), .A2(n699), .ZN(n742) );
  INV_X1 U569 ( .A(KEYINPUT95), .ZN(n759) );
  INV_X1 U570 ( .A(KEYINPUT64), .ZN(n766) );
  INV_X1 U571 ( .A(n956), .ZN(n778) );
  NAND2_X1 U572 ( .A1(n645), .A2(G81), .ZN(n571) );
  INV_X1 U573 ( .A(n836), .ZN(n825) );
  INV_X1 U574 ( .A(KEYINPUT13), .ZN(n574) );
  INV_X1 U575 ( .A(KEYINPUT73), .ZN(n585) );
  XNOR2_X1 U576 ( .A(n575), .B(n574), .ZN(n576) );
  NOR2_X1 U577 ( .A1(n577), .A2(n576), .ZN(n578) );
  INV_X1 U578 ( .A(KEYINPUT65), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n541), .A2(n540), .ZN(n542) );
  INV_X1 U580 ( .A(KEYINPUT100), .ZN(n828) );
  NOR2_X1 U581 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n630) );
  BUF_X1 U583 ( .A(n702), .Z(n970) );
  XNOR2_X1 U584 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n645), .A2(G89), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT4), .ZN(n525) );
  INV_X1 U588 ( .A(G651), .ZN(n527) );
  NOR2_X1 U589 ( .A1(n630), .A2(n527), .ZN(n649) );
  NAND2_X1 U590 ( .A1(G76), .A2(n649), .ZN(n524) );
  NAND2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(KEYINPUT5), .ZN(n534) );
  XOR2_X2 U593 ( .A(KEYINPUT1), .B(n528), .Z(n646) );
  NAND2_X1 U594 ( .A1(G63), .A2(n646), .ZN(n531) );
  NOR2_X1 U595 ( .A1(G651), .A2(n630), .ZN(n529) );
  XNOR2_X2 U596 ( .A(KEYINPUT66), .B(n529), .ZN(n653) );
  NAND2_X1 U597 ( .A1(G51), .A2(n653), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X4 U601 ( .A1(n541), .A2(n540), .ZN(n897) );
  NAND2_X1 U602 ( .A1(G114), .A2(n897), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT84), .ZN(n539) );
  NOR2_X1 U604 ( .A1(G2104), .A2(n540), .ZN(n691) );
  NAND2_X1 U605 ( .A1(G126), .A2(n691), .ZN(n537) );
  XOR2_X1 U606 ( .A(KEYINPUT83), .B(n537), .Z(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n548) );
  INV_X4 U608 ( .A(G2104), .ZN(n541) );
  XNOR2_X2 U609 ( .A(n542), .B(KEYINPUT17), .ZN(n690) );
  NAND2_X1 U610 ( .A1(G138), .A2(n690), .ZN(n544) );
  NOR2_X4 U611 ( .A1(G2105), .A2(n541), .ZN(n902) );
  NAND2_X1 U612 ( .A1(G102), .A2(n902), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n546) );
  INV_X1 U614 ( .A(KEYINPUT85), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n547) );
  NOR2_X2 U616 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U617 ( .A1(G64), .A2(n646), .ZN(n550) );
  NAND2_X1 U618 ( .A1(G52), .A2(n653), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G90), .A2(n645), .ZN(n552) );
  NAND2_X1 U621 ( .A1(G77), .A2(n649), .ZN(n551) );
  NAND2_X1 U622 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(KEYINPUT68), .B(n556), .ZN(G171) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  XOR2_X1 U627 ( .A(G2446), .B(G2451), .Z(n558) );
  XNOR2_X1 U628 ( .A(G2454), .B(KEYINPUT103), .ZN(n557) );
  XNOR2_X1 U629 ( .A(n558), .B(n557), .ZN(n565) );
  XOR2_X1 U630 ( .A(G2438), .B(G2430), .Z(n560) );
  XNOR2_X1 U631 ( .A(G2435), .B(G2443), .ZN(n559) );
  XNOR2_X1 U632 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U633 ( .A(n561), .B(G2427), .Z(n563) );
  XNOR2_X1 U634 ( .A(G1348), .B(G1341), .ZN(n562) );
  XNOR2_X1 U635 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U636 ( .A(n565), .B(n564), .ZN(n566) );
  AND2_X1 U637 ( .A1(n566), .A2(G14), .ZN(G401) );
  AND2_X1 U638 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U639 ( .A(G132), .ZN(G219) );
  INV_X1 U640 ( .A(G82), .ZN(G220) );
  INV_X1 U641 ( .A(G69), .ZN(G235) );
  INV_X1 U642 ( .A(G108), .ZN(G238) );
  INV_X1 U643 ( .A(G120), .ZN(G236) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U646 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n845) );
  NAND2_X1 U648 ( .A1(n845), .A2(G567), .ZN(n568) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U650 ( .A1(G56), .A2(n646), .ZN(n569) );
  XNOR2_X1 U651 ( .A(n569), .B(KEYINPUT71), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n570), .B(KEYINPUT14), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U654 ( .A1(G68), .A2(n649), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n578), .B(KEYINPUT72), .ZN(n580) );
  NAND2_X1 U657 ( .A1(G43), .A2(n653), .ZN(n579) );
  INV_X1 U658 ( .A(G860), .ZN(n602) );
  OR2_X1 U659 ( .A1(n970), .A2(n602), .ZN(G153) );
  NAND2_X1 U660 ( .A1(G301), .A2(G868), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G79), .A2(n649), .ZN(n582) );
  NAND2_X1 U662 ( .A1(G54), .A2(n653), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G66), .A2(n646), .ZN(n584) );
  NAND2_X1 U665 ( .A1(G92), .A2(n645), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U667 ( .A(n586), .B(n585), .ZN(n587) );
  NOR2_X1 U668 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X2 U669 ( .A(KEYINPUT15), .B(n589), .Z(n951) );
  OR2_X1 U670 ( .A1(n951), .A2(G868), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G65), .A2(n646), .ZN(n593) );
  NAND2_X1 U673 ( .A1(G53), .A2(n653), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G91), .A2(n645), .ZN(n595) );
  NAND2_X1 U676 ( .A1(G78), .A2(n649), .ZN(n594) );
  NAND2_X1 U677 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U678 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n598), .B(KEYINPUT69), .ZN(G299) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n599) );
  XNOR2_X1 U681 ( .A(n599), .B(KEYINPUT74), .ZN(n601) );
  INV_X1 U682 ( .A(G868), .ZN(n666) );
  NOR2_X1 U683 ( .A1(n666), .A2(G286), .ZN(n600) );
  NOR2_X1 U684 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n603), .A2(n951), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n970), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G868), .A2(n951), .ZN(n605) );
  NOR2_X1 U690 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U692 ( .A(KEYINPUT75), .B(n608), .Z(G282) );
  BUF_X1 U693 ( .A(n691), .Z(n898) );
  NAND2_X1 U694 ( .A1(G123), .A2(n898), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n902), .A2(G99), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G135), .A2(n612), .ZN(n614) );
  NAND2_X1 U699 ( .A1(G111), .A2(n897), .ZN(n613) );
  NAND2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n981) );
  XNOR2_X1 U702 ( .A(G2096), .B(n981), .ZN(n618) );
  INV_X1 U703 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G559), .A2(n951), .ZN(n619) );
  XNOR2_X1 U706 ( .A(n970), .B(n619), .ZN(n663) );
  NOR2_X1 U707 ( .A1(n663), .A2(G860), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G67), .A2(n646), .ZN(n621) );
  NAND2_X1 U709 ( .A1(G55), .A2(n653), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G93), .A2(n645), .ZN(n623) );
  NAND2_X1 U712 ( .A1(G80), .A2(n649), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U714 ( .A1(n625), .A2(n624), .ZN(n665) );
  XNOR2_X1 U715 ( .A(n626), .B(n665), .ZN(G145) );
  NAND2_X1 U716 ( .A1(G651), .A2(G74), .ZN(n628) );
  NAND2_X1 U717 ( .A1(G49), .A2(n653), .ZN(n627) );
  NAND2_X1 U718 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U719 ( .A1(n646), .A2(n629), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G88), .A2(n645), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G75), .A2(n649), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U725 ( .A1(G62), .A2(n646), .ZN(n636) );
  NAND2_X1 U726 ( .A1(G50), .A2(n653), .ZN(n635) );
  NAND2_X1 U727 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U728 ( .A1(n638), .A2(n637), .ZN(G166) );
  AND2_X1 U729 ( .A1(n646), .A2(G60), .ZN(n642) );
  NAND2_X1 U730 ( .A1(G85), .A2(n645), .ZN(n640) );
  NAND2_X1 U731 ( .A1(G72), .A2(n649), .ZN(n639) );
  NAND2_X1 U732 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U733 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U734 ( .A1(G47), .A2(n653), .ZN(n643) );
  NAND2_X1 U735 ( .A1(n644), .A2(n643), .ZN(G290) );
  NAND2_X1 U736 ( .A1(G86), .A2(n645), .ZN(n648) );
  NAND2_X1 U737 ( .A1(G61), .A2(n646), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G48), .A2(n653), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(G305) );
  XNOR2_X1 U744 ( .A(KEYINPUT19), .B(KEYINPUT76), .ZN(n657) );
  XNOR2_X1 U745 ( .A(G288), .B(KEYINPUT77), .ZN(n656) );
  XNOR2_X1 U746 ( .A(n657), .B(n656), .ZN(n660) );
  XNOR2_X1 U747 ( .A(G166), .B(G290), .ZN(n658) );
  XNOR2_X1 U748 ( .A(n658), .B(G299), .ZN(n659) );
  XNOR2_X1 U749 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U750 ( .A(G305), .B(n665), .ZN(n661) );
  XNOR2_X1 U751 ( .A(n662), .B(n661), .ZN(n851) );
  XOR2_X1 U752 ( .A(n663), .B(n851), .Z(n664) );
  NAND2_X1 U753 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U756 ( .A(KEYINPUT78), .B(n669), .Z(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XNOR2_X1 U758 ( .A(n670), .B(KEYINPUT79), .ZN(n671) );
  XNOR2_X1 U759 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XOR2_X1 U763 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U765 ( .A1(G236), .A2(G238), .ZN(n676) );
  NOR2_X1 U766 ( .A1(G235), .A2(G237), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U768 ( .A(KEYINPUT80), .B(n677), .ZN(n850) );
  NAND2_X1 U769 ( .A1(n850), .A2(G567), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U772 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G96), .A2(n680), .ZN(n849) );
  NAND2_X1 U774 ( .A1(G2106), .A2(n849), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U776 ( .A(KEYINPUT81), .B(n683), .ZN(G319) );
  INV_X1 U777 ( .A(G319), .ZN(n919) );
  NAND2_X1 U778 ( .A1(G661), .A2(G483), .ZN(n684) );
  XNOR2_X1 U779 ( .A(KEYINPUT82), .B(n684), .ZN(n685) );
  NOR2_X1 U780 ( .A1(n919), .A2(n685), .ZN(n848) );
  NAND2_X1 U781 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(G101), .A2(n902), .ZN(n686) );
  XOR2_X1 U783 ( .A(KEYINPUT23), .B(n686), .Z(n689) );
  NAND2_X1 U784 ( .A1(G113), .A2(n897), .ZN(n687) );
  XOR2_X1 U785 ( .A(KEYINPUT67), .B(n687), .Z(n688) );
  NAND2_X1 U786 ( .A1(n689), .A2(n688), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G137), .A2(n690), .ZN(n693) );
  NAND2_X1 U788 ( .A1(G125), .A2(n691), .ZN(n692) );
  NAND2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n695) );
  NOR2_X1 U790 ( .A1(n697), .A2(n695), .ZN(G160) );
  INV_X1 U791 ( .A(G166), .ZN(G303) );
  NOR2_X2 U792 ( .A1(G164), .A2(G1384), .ZN(n795) );
  INV_X1 U793 ( .A(G40), .ZN(n694) );
  OR2_X1 U794 ( .A1(n695), .A2(n694), .ZN(n696) );
  INV_X1 U795 ( .A(n794), .ZN(n699) );
  AND2_X2 U796 ( .A1(n795), .A2(n699), .ZN(n724) );
  XOR2_X1 U797 ( .A(n698), .B(KEYINPUT26), .Z(n701) );
  NAND2_X1 U798 ( .A1(n742), .A2(G1341), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U801 ( .A1(n706), .A2(n951), .ZN(n705) );
  XNOR2_X1 U802 ( .A(n705), .B(n704), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n706), .A2(n951), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n724), .A2(G1348), .ZN(n708) );
  NOR2_X1 U805 ( .A1(G2067), .A2(n742), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n717) );
  INV_X1 U809 ( .A(G299), .ZN(n958) );
  NAND2_X1 U810 ( .A1(n724), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U811 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  XNOR2_X1 U812 ( .A(KEYINPUT89), .B(G1956), .ZN(n932) );
  NOR2_X1 U813 ( .A1(n932), .A2(n724), .ZN(n714) );
  NOR2_X1 U814 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n958), .A2(n718), .ZN(n716) );
  NAND2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U817 ( .A1(n958), .A2(n718), .ZN(n719) );
  XOR2_X1 U818 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U819 ( .A1(n721), .A2(n720), .ZN(n723) );
  INV_X1 U820 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U821 ( .A(n723), .B(n722), .ZN(n727) );
  NAND2_X1 U822 ( .A1(G1961), .A2(n742), .ZN(n726) );
  XOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .Z(n1017) );
  NAND2_X1 U824 ( .A1(n724), .A2(n1017), .ZN(n725) );
  NAND2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n727), .A2(n516), .ZN(n740) );
  NAND2_X1 U827 ( .A1(G301), .A2(n728), .ZN(n729) );
  XOR2_X1 U828 ( .A(KEYINPUT92), .B(n729), .Z(n736) );
  NAND2_X1 U829 ( .A1(G8), .A2(n742), .ZN(n741) );
  NOR2_X1 U830 ( .A1(G2084), .A2(n742), .ZN(n751) );
  NOR2_X1 U831 ( .A1(n754), .A2(n751), .ZN(n730) );
  NAND2_X1 U832 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U833 ( .A(n731), .B(KEYINPUT30), .ZN(n732) );
  NOR2_X1 U834 ( .A1(n732), .A2(G168), .ZN(n734) );
  NOR2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U836 ( .A1(n740), .A2(n520), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n752), .A2(G286), .ZN(n749) );
  INV_X1 U838 ( .A(G8), .ZN(n747) );
  INV_X1 U839 ( .A(n741), .ZN(n763) );
  INV_X1 U840 ( .A(n763), .ZN(n787) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n787), .ZN(n744) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n742), .ZN(n743) );
  NOR2_X1 U843 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n745), .A2(G303), .ZN(n746) );
  OR2_X1 U845 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U846 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U847 ( .A(n750), .B(n519), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n751), .A2(G8), .ZN(n756) );
  INV_X1 U849 ( .A(n752), .ZN(n753) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U852 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U853 ( .A(n760), .B(n759), .ZN(n785) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n773) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U856 ( .A1(n773), .A2(n761), .ZN(n965) );
  XNOR2_X1 U857 ( .A(KEYINPUT96), .B(n965), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n785), .A2(n762), .ZN(n765) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n961) );
  AND2_X1 U860 ( .A1(n763), .A2(n961), .ZN(n764) );
  NAND2_X1 U861 ( .A1(n765), .A2(n764), .ZN(n767) );
  XNOR2_X1 U862 ( .A(n767), .B(n766), .ZN(n768) );
  INV_X1 U863 ( .A(KEYINPUT97), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n768), .A2(n517), .ZN(n770) );
  INV_X1 U865 ( .A(KEYINPUT33), .ZN(n769) );
  NAND2_X1 U866 ( .A1(n770), .A2(n769), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n773), .A2(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U868 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n773), .A2(KEYINPUT97), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U871 ( .A1(n787), .A2(n776), .ZN(n779) );
  XOR2_X1 U872 ( .A(G1981), .B(KEYINPUT98), .Z(n777) );
  XNOR2_X1 U873 ( .A(G305), .B(n777), .ZN(n956) );
  NOR2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n792) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U877 ( .A(n782), .B(KEYINPUT24), .Z(n783) );
  OR2_X1 U878 ( .A1(n787), .A2(n783), .ZN(n790) );
  NOR2_X1 U879 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U880 ( .A1(G8), .A2(n784), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n789) );
  AND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U884 ( .A(n793), .B(KEYINPUT99), .ZN(n827) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n840) );
  INV_X1 U886 ( .A(n840), .ZN(n815) );
  XNOR2_X1 U887 ( .A(G1986), .B(G290), .ZN(n967) );
  NAND2_X1 U888 ( .A1(G107), .A2(n897), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G119), .A2(n898), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G131), .A2(n612), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G95), .A2(n902), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U894 ( .A(KEYINPUT86), .B(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(n803), .B(KEYINPUT87), .ZN(n917) );
  NAND2_X1 U897 ( .A1(G1991), .A2(n917), .ZN(n813) );
  NAND2_X1 U898 ( .A1(G141), .A2(n612), .ZN(n804) );
  XNOR2_X1 U899 ( .A(n804), .B(KEYINPUT88), .ZN(n811) );
  NAND2_X1 U900 ( .A1(G117), .A2(n897), .ZN(n806) );
  NAND2_X1 U901 ( .A1(G129), .A2(n898), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n902), .A2(G105), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT38), .B(n807), .Z(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n911) );
  NAND2_X1 U907 ( .A1(G1996), .A2(n911), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n993) );
  NOR2_X1 U909 ( .A1(n967), .A2(n993), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n826) );
  XNOR2_X1 U911 ( .A(KEYINPUT37), .B(G2067), .ZN(n838) );
  NAND2_X1 U912 ( .A1(G140), .A2(n612), .ZN(n817) );
  NAND2_X1 U913 ( .A1(G104), .A2(n902), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U915 ( .A(KEYINPUT34), .B(n818), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G116), .A2(n897), .ZN(n820) );
  NAND2_X1 U917 ( .A1(G128), .A2(n898), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U919 ( .A(KEYINPUT35), .B(n821), .Z(n822) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT36), .B(n824), .ZN(n914) );
  NOR2_X1 U922 ( .A1(n838), .A2(n914), .ZN(n983) );
  NAND2_X1 U923 ( .A1(n840), .A2(n983), .ZN(n836) );
  AND2_X1 U924 ( .A1(n827), .A2(n518), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n843) );
  NOR2_X1 U926 ( .A1(G1996), .A2(n911), .ZN(n988) );
  NOR2_X1 U927 ( .A1(G1991), .A2(n917), .ZN(n982) );
  NOR2_X1 U928 ( .A1(G1986), .A2(G290), .ZN(n830) );
  XOR2_X1 U929 ( .A(n830), .B(KEYINPUT101), .Z(n831) );
  NOR2_X1 U930 ( .A1(n982), .A2(n831), .ZN(n832) );
  NOR2_X1 U931 ( .A1(n832), .A2(n993), .ZN(n833) );
  NOR2_X1 U932 ( .A1(n988), .A2(n833), .ZN(n834) );
  XNOR2_X1 U933 ( .A(KEYINPUT39), .B(n834), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n835), .B(KEYINPUT102), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n838), .A2(n914), .ZN(n995) );
  NAND2_X1 U937 ( .A1(n839), .A2(n995), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n844), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  NOR2_X1 U948 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(n970), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(G301), .B(n951), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n854), .B(G286), .ZN(n855) );
  NOR2_X1 U954 ( .A1(G37), .A2(n855), .ZN(G397) );
  XOR2_X1 U955 ( .A(G1981), .B(G1966), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1961), .B(G1956), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n867) );
  XOR2_X1 U958 ( .A(G2474), .B(KEYINPUT107), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1996), .B(KEYINPUT41), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(G1976), .B(G1971), .Z(n861) );
  XNOR2_X1 U962 ( .A(G1991), .B(G1986), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(G229) );
  XOR2_X1 U968 ( .A(G2096), .B(KEYINPUT43), .Z(n869) );
  XNOR2_X1 U969 ( .A(G2072), .B(G2678), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(n870), .B(KEYINPUT104), .Z(n872) );
  XNOR2_X1 U972 ( .A(G2067), .B(G2090), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT42), .B(G2100), .Z(n874) );
  XNOR2_X1 U975 ( .A(G2078), .B(G2084), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(G227) );
  NAND2_X1 U978 ( .A1(G100), .A2(n902), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G112), .A2(n897), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G124), .A2(n898), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G136), .A2(n612), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n880), .B(KEYINPUT108), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n886) );
  XNOR2_X1 U988 ( .A(n981), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G118), .A2(n897), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G130), .A2(n898), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G142), .A2(n612), .ZN(n890) );
  NAND2_X1 U994 ( .A1(G106), .A2(n902), .ZN(n889) );
  NAND2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U996 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  XNOR2_X1 U997 ( .A(KEYINPUT109), .B(n892), .ZN(n893) );
  NOR2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U999 ( .A(n896), .B(n895), .Z(n909) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n897), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n898), .ZN(n899) );
  NAND2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n901), .B(KEYINPUT47), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n902), .ZN(n903) );
  NAND2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n612), .A2(G139), .ZN(n905) );
  XOR2_X1 U1007 ( .A(KEYINPUT110), .B(n905), .Z(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n997) );
  XNOR2_X1 U1009 ( .A(n997), .B(G162), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(G164), .B(G160), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1014 ( .A(n915), .B(n914), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n919), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(G397), .A2(n921), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n924), .A2(G395), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1024 ( .A(G308), .ZN(G225) );
  XOR2_X1 U1025 ( .A(G1976), .B(G23), .Z(n928) );
  XNOR2_X1 U1026 ( .A(G1986), .B(KEYINPUT127), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n926), .B(G24), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(G22), .B(G1971), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT58), .B(n931), .Z(n948) );
  XOR2_X1 U1032 ( .A(G1961), .B(G5), .Z(n942) );
  XNOR2_X1 U1033 ( .A(G20), .B(n932), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(G6), .B(G1981), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1038 ( .A(KEYINPUT59), .B(G1348), .Z(n937) );
  XNOR2_X1 U1039 ( .A(G4), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(KEYINPUT60), .B(n940), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1043 ( .A(G21), .B(G1966), .Z(n943) );
  XNOR2_X1 U1044 ( .A(KEYINPUT125), .B(n943), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1046 ( .A(KEYINPUT126), .B(n946), .Z(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1048 ( .A(KEYINPUT61), .B(n949), .Z(n950) );
  NOR2_X1 U1049 ( .A1(G16), .A2(n950), .ZN(n979) );
  XNOR2_X1 U1050 ( .A(KEYINPUT56), .B(G16), .ZN(n976) );
  XOR2_X1 U1051 ( .A(G1348), .B(n951), .Z(n953) );
  XNOR2_X1 U1052 ( .A(G301), .B(G1961), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n974) );
  XNOR2_X1 U1054 ( .A(G168), .B(G1966), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(n954), .B(KEYINPUT122), .ZN(n955) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(n957), .B(KEYINPUT57), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(n958), .B(G1956), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(KEYINPUT123), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n970), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1070 ( .A(KEYINPUT124), .B(n977), .Z(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n1008) );
  XOR2_X1 U1072 ( .A(G2084), .B(G160), .Z(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n985) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT113), .B(n986), .ZN(n991) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT51), .B(n989), .Z(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n994), .B(KEYINPUT114), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(G2072), .B(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G164), .B(G2078), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT115), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT50), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1004), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1028) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1028), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(G29), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  XNOR2_X1 U1095 ( .A(KEYINPUT54), .B(G34), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT119), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G2084), .B(n1010), .ZN(n1027) );
  XNOR2_X1 U1098 ( .A(G2090), .B(G35), .ZN(n1025) );
  XOR2_X1 U1099 ( .A(G1991), .B(G25), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(G28), .A2(n1011), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT117), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G2067), .B(G26), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(G33), .B(G2072), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G1996), .B(G32), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1017), .B(G27), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(KEYINPUT118), .B(n1020), .Z(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(KEYINPUT53), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(n1028), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(G29), .B(KEYINPUT120), .Z(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(G11), .ZN(n1033) );
  XOR2_X1 U1118 ( .A(KEYINPUT121), .B(n1033), .Z(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

