//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(new_n212), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT2), .B(G226), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  OR2_X1    g0040(.A1(KEYINPUT5), .A2(G41), .ZN(new_n241));
  NAND2_X1  g0041(.A1(KEYINPUT5), .A2(G41), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(new_n244), .A3(G45), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT65), .B1(new_n247), .B2(new_n210), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT65), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n211), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n245), .A2(G270), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n244), .A2(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n241), .B2(new_n242), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(new_n248), .A3(G274), .A4(new_n250), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G116), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(new_n210), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n244), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(G116), .A3(new_n256), .A4(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n210), .B1(G20), .B2(new_n258), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G283), .ZN(new_n265));
  INV_X1    g0065(.A(G20), .ZN(new_n266));
  INV_X1    g0066(.A(G97), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n265), .B(new_n266), .C1(G33), .C2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n264), .A2(KEYINPUT20), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT20), .B1(new_n264), .B2(new_n268), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n259), .B(new_n263), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  OAI211_X1 g0075(.A(G257), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G303), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n247), .A2(new_n210), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n255), .A2(G179), .A3(new_n271), .A4(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n251), .A3(new_n254), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(KEYINPUT21), .A3(new_n271), .A4(G169), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G169), .A3(new_n271), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT21), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n271), .B1(new_n286), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n288), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G116), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n266), .B2(G107), .ZN(new_n300));
  INV_X1    g0100(.A(G107), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(KEYINPUT23), .A3(G20), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n266), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT22), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(KEYINPUT86), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n304), .A2(new_n306), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT24), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n303), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n260), .A2(new_n210), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n261), .A2(new_n256), .A3(new_n262), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT25), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n256), .B2(G107), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n256), .A2(new_n317), .A3(G107), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n316), .A2(new_n301), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(G257), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n323));
  OAI211_X1 g0123(.A(G250), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n324));
  INV_X1    g0124(.A(G294), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n323), .B(new_n324), .C1(new_n278), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n283), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n245), .A2(G264), .A3(new_n248), .A4(new_n250), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n254), .A3(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(new_n293), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(G200), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n315), .A2(new_n322), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n327), .A2(new_n328), .A3(new_n333), .A4(new_n254), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n261), .B1(new_n310), .B2(new_n312), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n334), .B(new_n336), .C1(new_n337), .C2(new_n321), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n296), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n266), .A3(new_n278), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT68), .B1(G20), .B2(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G50), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT67), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n278), .B2(G20), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n266), .A2(KEYINPUT67), .A3(G33), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n348), .B1(new_n266), .B2(G68), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT11), .A3(new_n314), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n314), .B1(new_n244), .B2(G20), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n256), .A2(KEYINPUT12), .A3(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT12), .B1(new_n256), .B2(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(G68), .A2(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n354), .B2(new_n314), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n275), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n225), .A2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(new_n272), .C2(new_n273), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n368), .A2(KEYINPUT70), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT70), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(new_n283), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G41), .ZN(new_n374));
  INV_X1    g0174(.A(G45), .ZN(new_n375));
  AOI21_X1  g0175(.A(G1), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n248), .A2(new_n377), .A3(new_n250), .A4(G238), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n248), .A2(new_n250), .A3(G274), .A4(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT13), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n368), .A2(new_n369), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT70), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n368), .A2(KEYINPUT70), .A3(new_n369), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n283), .ZN(new_n386));
  INV_X1    g0186(.A(new_n380), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n381), .A2(G179), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n381), .A2(new_n392), .A3(G179), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n373), .A2(KEYINPUT13), .A3(new_n380), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n388), .B1(new_n386), .B2(new_n387), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n381), .A2(new_n389), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(G169), .ZN(new_n401));
  AND4_X1   g0201(.A1(new_n364), .A2(new_n394), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n400), .B1(new_n399), .B2(G169), .ZN(new_n403));
  AOI211_X1 g0203(.A(KEYINPUT14), .B(new_n335), .C1(new_n381), .C2(new_n389), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n364), .B1(new_n405), .B2(new_n394), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n363), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n248), .A2(new_n377), .A3(new_n250), .A4(G232), .ZN(new_n409));
  NOR2_X1   g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n365), .B2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n279), .A2(new_n280), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(G33), .B2(G87), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n409), .B(new_n379), .C1(new_n413), .C2(new_n372), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT75), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n283), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT75), .B1(new_n413), .B2(new_n372), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n409), .A2(new_n379), .A3(new_n293), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n416), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT8), .B(G58), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT66), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G58), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n356), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n256), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n279), .A2(new_n266), .A3(new_n280), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT7), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n266), .A4(new_n280), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(KEYINPUT74), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(G68), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(G58), .B(G68), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n345), .A2(G159), .B1(new_n443), .B2(G20), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT16), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n272), .A2(new_n273), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT7), .B1(new_n446), .B2(new_n266), .ZN(new_n447));
  INV_X1    g0247(.A(new_n438), .ZN(new_n448));
  OAI21_X1  g0248(.A(G68), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT16), .A3(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n314), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n425), .B(new_n434), .C1(new_n445), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n408), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n434), .B1(new_n445), .B2(new_n451), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n421), .A2(new_n422), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n379), .A2(new_n409), .A3(new_n333), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(new_n457), .B1(new_n414), .B2(new_n335), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT18), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n442), .A2(new_n444), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G68), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n437), .B2(new_n438), .ZN(new_n465));
  INV_X1    g0265(.A(new_n444), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n261), .B1(new_n467), .B2(KEYINPUT16), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n433), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n425), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n455), .A2(new_n458), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n454), .A2(new_n460), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n399), .A2(G200), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n381), .A2(G190), .A3(new_n389), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n362), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n431), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n351), .A2(new_n352), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n345), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n261), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n256), .A2(G50), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n356), .B2(G50), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n412), .A2(G223), .A3(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n412), .A2(G222), .A3(new_n275), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n349), .C2(new_n412), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n283), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n248), .A2(new_n377), .A3(new_n250), .A4(G226), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(new_n379), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n333), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n492), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n335), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n257), .A2(new_n349), .ZN(new_n498));
  INV_X1    g0298(.A(new_n356), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n349), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT15), .B(G87), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n479), .B1(G20), .B2(G77), .ZN(new_n503));
  INV_X1    g0303(.A(new_n345), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n426), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n500), .B1(new_n505), .B2(new_n314), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G232), .A2(G1698), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n275), .A2(G238), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n412), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n283), .C1(G107), .C2(new_n412), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n248), .A2(new_n377), .A3(new_n250), .A4(G244), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n379), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n333), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n335), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(G200), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n506), .C1(new_n293), .C2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n494), .A2(new_n293), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n415), .B1(new_n490), .B2(new_n492), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT9), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n483), .B2(new_n485), .ZN(new_n525));
  INV_X1    g0325(.A(new_n485), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n482), .A2(KEYINPUT9), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT10), .B1(new_n522), .B2(KEYINPUT69), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n523), .B(new_n529), .C1(new_n525), .C2(new_n527), .ZN(new_n532));
  AOI211_X1 g0332(.A(new_n497), .B(new_n520), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AND4_X1   g0333(.A1(new_n407), .A2(new_n474), .A3(new_n477), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n502), .A2(new_n256), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n266), .B(G68), .C1(new_n272), .C2(new_n273), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n267), .B1(new_n351), .B2(new_n352), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n266), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n267), .A3(new_n301), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n540), .B2(new_n543), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n537), .B1(new_n538), .B2(KEYINPUT19), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n261), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT82), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n353), .B2(new_n267), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT83), .A4(new_n537), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n536), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n316), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G87), .ZN(new_n558));
  OAI211_X1 g0358(.A(G244), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n559));
  OAI211_X1 g0359(.A(G238), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n297), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n283), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n252), .A2(G274), .ZN(new_n563));
  INV_X1    g0363(.A(G250), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n252), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(new_n248), .A3(new_n250), .A4(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n562), .A2(KEYINPUT81), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT81), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(KEYINPUT81), .A3(new_n566), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(G190), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n556), .A2(new_n558), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n544), .A2(new_n545), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n537), .B1(new_n538), .B2(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n547), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n555), .A3(new_n314), .ZN(new_n579));
  INV_X1    g0379(.A(new_n536), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n316), .A2(new_n501), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT84), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n335), .B1(new_n567), .B2(new_n568), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n572), .A2(new_n333), .A3(new_n573), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n575), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n245), .A2(G257), .A3(new_n248), .A4(new_n250), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n254), .ZN(new_n590));
  OAI211_X1 g0390(.A(G244), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n591), .A2(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(KEYINPUT78), .A3(new_n592), .ZN(new_n597));
  OAI211_X1 g0397(.A(G250), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n598), .A2(new_n265), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n590), .B1(new_n600), .B2(new_n283), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n439), .A2(G107), .A3(new_n441), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  AND2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G97), .A2(G107), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n301), .A2(KEYINPUT6), .A3(G97), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n266), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n344), .ZN(new_n610));
  NOR3_X1   g0410(.A1(KEYINPUT68), .A2(G20), .A3(G33), .ZN(new_n611));
  OAI21_X1  g0411(.A(G77), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT77), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n345), .A2(new_n614), .A3(G77), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n261), .B1(new_n603), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n256), .A2(G97), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n557), .B2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(G200), .B1(new_n601), .B2(KEYINPUT79), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT79), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n623), .B(new_n590), .C1(new_n600), .C2(new_n283), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n602), .B(new_n621), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n589), .A2(new_n254), .ZN(new_n626));
  INV_X1    g0426(.A(new_n597), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n598), .B(new_n265), .C1(new_n591), .C2(new_n592), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT78), .B1(new_n591), .B2(new_n592), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(G179), .B(new_n626), .C1(new_n630), .C2(new_n372), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n335), .B2(new_n601), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT80), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n603), .A2(new_n616), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n314), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n619), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n617), .A2(KEYINPUT80), .A3(new_n620), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n587), .A2(new_n588), .A3(new_n625), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n625), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n575), .A2(new_n586), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT85), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n341), .B(new_n535), .C1(new_n639), .C2(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n531), .A2(new_n532), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n454), .A2(new_n470), .ZN(new_n645));
  INV_X1    g0445(.A(new_n517), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n477), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n407), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n460), .A2(new_n472), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n644), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(new_n496), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n336), .A2(new_n334), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n315), .B2(new_n322), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n291), .A2(new_n285), .A3(new_n287), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT87), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n338), .A2(new_n657), .A3(new_n291), .A4(new_n288), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n570), .A2(G200), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n556), .A2(new_n558), .A3(new_n574), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n570), .A2(new_n335), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n583), .A2(new_n585), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n332), .A3(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n659), .A2(new_n640), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT26), .B1(new_n641), .B2(new_n638), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n663), .B(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n626), .B1(new_n630), .B2(new_n372), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G169), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n621), .B1(new_n670), .B2(new_n631), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n661), .A3(new_n663), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n666), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n534), .B1(new_n665), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n652), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n244), .A2(new_n266), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n271), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g0483(.A(new_n655), .B(new_n295), .S(new_n683), .Z(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n682), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n315), .B2(new_n322), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n339), .A2(new_n687), .B1(new_n338), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n655), .A2(new_n686), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n339), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n654), .B2(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n543), .A2(G116), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT89), .ZN(new_n695));
  INV_X1    g0495(.A(new_n207), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n244), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n214), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT28), .Z(new_n701));
  NAND4_X1  g0501(.A1(new_n295), .A2(new_n338), .A3(new_n332), .A4(new_n686), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n642), .B2(new_n639), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n286), .A2(new_n333), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n327), .A2(new_n328), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n601), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n572), .A2(new_n573), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n709), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n706), .A2(new_n286), .A3(new_n333), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT30), .A4(new_n601), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n286), .A2(new_n333), .A3(new_n570), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n669), .A3(new_n329), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n682), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n725), .B(new_n686), .C1(new_n665), .C2(new_n674), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n672), .B1(new_n641), .B2(new_n638), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n671), .A2(new_n661), .A3(new_n663), .A4(KEYINPUT26), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n669), .A2(new_n623), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G200), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n602), .A2(new_n621), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n635), .A2(new_n633), .A3(new_n619), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT80), .B1(new_n617), .B2(new_n620), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n737), .B2(new_n632), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n661), .A2(new_n663), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n338), .A2(new_n291), .A3(new_n288), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n332), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n730), .A2(new_n741), .A3(new_n668), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n725), .B1(new_n742), .B2(new_n686), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n724), .A2(new_n727), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n701), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(G13), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n244), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n685), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n684), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n696), .A2(new_n446), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G355), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G116), .B2(new_n207), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n236), .A2(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n696), .A2(new_n412), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n375), .B2(new_n699), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n210), .B1(G20), .B2(new_n335), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT90), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT90), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n750), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n764), .ZN(new_n771));
  NAND2_X1  g0571(.A1(G20), .A2(G179), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n266), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n266), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n779), .B1(new_n325), .B2(new_n781), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n412), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n773), .A2(new_n786), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n772), .A2(new_n293), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(new_n790), .B2(new_n791), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n774), .A2(new_n293), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G326), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n783), .A2(new_n293), .A3(G200), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n785), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  INV_X1    g0602(.A(new_n775), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n464), .ZN(new_n804));
  INV_X1    g0604(.A(new_n796), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(G159), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n202), .B1(new_n806), .B2(KEYINPUT32), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(KEYINPUT32), .C2(new_n806), .ZN(new_n808));
  INV_X1    g0608(.A(new_n784), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G87), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n301), .B2(new_n799), .ZN(new_n811));
  INV_X1    g0611(.A(new_n781), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n446), .B(new_n811), .C1(G97), .C2(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n794), .A2(new_n429), .B1(new_n791), .B2(new_n349), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT91), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n808), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n802), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT93), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n771), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(KEYINPUT93), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n770), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n767), .B(KEYINPUT94), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n684), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n752), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  OAI21_X1  g0626(.A(new_n686), .B1(new_n665), .B2(new_n674), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n517), .B(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n507), .A2(new_n682), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(new_n519), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n517), .A2(new_n686), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT97), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n686), .B(new_n834), .C1(new_n665), .C2(new_n674), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n724), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n750), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n724), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n764), .A2(new_n765), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n750), .B1(new_n844), .B2(G77), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n805), .A2(new_n782), .B1(new_n784), .B2(new_n301), .ZN(new_n846));
  INV_X1    g0646(.A(new_n799), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(G87), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n412), .B1(G294), .B2(new_n793), .ZN(new_n849));
  INV_X1    g0649(.A(new_n791), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G311), .A2(new_n788), .B1(new_n850), .B2(G116), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n812), .A2(G97), .B1(new_n775), .B2(G283), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT95), .B(G143), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n850), .A2(G159), .B1(new_n855), .B2(new_n793), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n803), .B2(new_n857), .C1(new_n858), .C2(new_n805), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n847), .A2(G68), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n446), .B1(new_n788), .B2(G132), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n812), .A2(G58), .B1(new_n809), .B2(G50), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n859), .A2(new_n860), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n853), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n845), .B1(new_n867), .B2(new_n764), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n834), .B2(new_n766), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n842), .A2(new_n869), .ZN(G384));
  OAI21_X1  g0670(.A(G77), .B1(new_n429), .B2(new_n464), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n214), .A2(new_n871), .B1(G50), .B2(new_n464), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G1), .A3(new_n746), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT98), .Z(new_n874));
  NAND2_X1  g0674(.A1(new_n607), .A2(new_n608), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n258), .B(new_n212), .C1(new_n875), .C2(KEYINPUT35), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(KEYINPUT35), .B2(new_n875), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT36), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  XNOR2_X1  g0680(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT100), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n680), .B(KEYINPUT99), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n469), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n455), .A2(KEYINPUT100), .A3(new_n883), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n459), .A2(new_n452), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n458), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n468), .B1(KEYINPUT16), .B2(new_n467), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n891), .A2(new_n680), .B1(new_n892), .B2(new_n434), .ZN(new_n893));
  INV_X1    g0693(.A(new_n452), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n680), .B1(new_n892), .B2(new_n434), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n473), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n363), .A2(new_n682), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n407), .A2(new_n477), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n391), .A2(new_n393), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n398), .A2(new_n401), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT73), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n405), .A2(new_n364), .A3(new_n394), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n477), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n363), .B(new_n682), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n642), .A2(new_n639), .ZN(new_n914));
  INV_X1    g0714(.A(new_n702), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n719), .A2(new_n720), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n835), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n903), .B1(new_n919), .B2(KEYINPUT102), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n834), .B1(new_n703), .B2(new_n721), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n905), .B2(new_n912), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n881), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n455), .A2(KEYINPUT100), .A3(new_n883), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT100), .B1(new_n455), .B2(new_n883), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n459), .A2(new_n452), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT37), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n890), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n473), .A2(new_n928), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT103), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT103), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n930), .A2(new_n890), .B1(new_n473), .B2(new_n928), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n902), .B(new_n936), .C1(new_n937), .C2(KEYINPUT38), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n913), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n925), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n535), .A2(new_n722), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n723), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n534), .B1(new_n727), .B2(new_n743), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n652), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n933), .B2(new_n934), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n902), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n407), .A2(new_n682), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n828), .A2(new_n682), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n837), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n901), .A2(new_n902), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(new_n913), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n650), .A2(new_n884), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n947), .B(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n945), .A2(new_n959), .B1(new_n244), .B2(new_n747), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT104), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n945), .A2(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(KEYINPUT104), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n880), .B1(new_n963), .B2(new_n964), .ZN(G367));
  OAI21_X1  g0765(.A(new_n768), .B1(new_n207), .B2(new_n501), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n231), .A2(new_n758), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n750), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n803), .A2(new_n325), .B1(new_n799), .B2(new_n267), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G311), .B2(new_n796), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n781), .A2(new_n301), .B1(new_n791), .B2(new_n798), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n412), .B1(new_n788), .B2(G317), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n784), .B2(new_n258), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n793), .A2(G303), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n799), .A2(new_n349), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G159), .B2(new_n775), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n429), .B2(new_n784), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n812), .A2(G68), .B1(new_n796), .B2(new_n855), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n446), .B1(new_n788), .B2(G137), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n850), .A2(G50), .B1(G150), .B2(new_n793), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n974), .A2(new_n980), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT47), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(new_n764), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n968), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n556), .A2(new_n558), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n682), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n739), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n668), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n993), .B1(new_n997), .B2(new_n823), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n738), .B1(new_n621), .B2(new_n686), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n671), .A2(new_n682), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n691), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT42), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n338), .B1(new_n999), .B2(new_n1000), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n638), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n686), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT105), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n997), .B(KEYINPUT43), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n689), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n1001), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1015), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1001), .A2(new_n692), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT45), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n1001), .A2(new_n692), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT44), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1016), .A2(KEYINPUT106), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n691), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n690), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n688), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n685), .B(new_n1028), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n744), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n697), .B(KEYINPUT41), .Z(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n749), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n998), .B1(new_n1018), .B2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(new_n1029), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(new_n744), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n744), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n697), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n688), .A2(new_n823), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n228), .A2(new_n375), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1040), .A2(new_n757), .B1(new_n695), .B2(new_n753), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(G50), .B2(new_n426), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n375), .C1(new_n464), .C2(new_n349), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(G50), .A3(new_n426), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1044), .A2(new_n695), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n301), .B2(new_n696), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n750), .B1(new_n1048), .B2(new_n769), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n794), .A2(new_n202), .B1(new_n791), .B2(new_n464), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n446), .B(new_n1050), .C1(G150), .C2(new_n788), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G159), .A2(new_n796), .B1(new_n847), .B2(G97), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n812), .A2(new_n502), .B1(new_n809), .B2(G77), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n478), .A2(new_n775), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n850), .A2(G303), .B1(G317), .B2(new_n793), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n803), .B2(new_n790), .C1(new_n792), .C2(new_n805), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n812), .A2(G283), .B1(new_n809), .B2(G294), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n412), .B1(new_n788), .B2(G326), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n258), .C2(new_n799), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1039), .B(new_n1049), .C1(new_n1068), .C2(new_n764), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1035), .B2(new_n749), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1038), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT110), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1038), .A2(KEYINPUT110), .A3(new_n1070), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(G393));
  NAND2_X1  g0875(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1020), .A2(new_n1022), .A3(new_n689), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n749), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n750), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n768), .B1(new_n267), .B2(new_n207), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n239), .B2(new_n757), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT111), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n781), .A2(new_n349), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n803), .A2(new_n202), .B1(new_n799), .B2(new_n542), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G68), .C2(new_n809), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n446), .B1(new_n788), .B2(new_n855), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n426), .C2(new_n791), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n796), .A2(G150), .B1(G159), .B2(new_n793), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n812), .A2(G116), .B1(G294), .B2(new_n850), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n782), .B2(new_n803), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT113), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n412), .B1(new_n788), .B2(G322), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n301), .B2(new_n799), .C1(new_n798), .C2(new_n784), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT112), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n796), .A2(G317), .B1(G311), .B2(new_n793), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1089), .A2(new_n1091), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1084), .B1(new_n764), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n767), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1001), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n697), .B1(new_n1025), .B2(new_n1037), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1108), .A2(new_n1037), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1078), .B(new_n1106), .C1(new_n1107), .C2(new_n1109), .ZN(G390));
  NAND2_X1  g0910(.A1(new_n949), .A2(new_n950), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n765), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n803), .A2(new_n301), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1085), .B(new_n1113), .C1(G283), .C2(new_n796), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n794), .A2(new_n258), .B1(new_n787), .B2(new_n325), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n412), .B(new_n1115), .C1(G97), .C2(new_n850), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n810), .A3(new_n862), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n791), .A2(new_n1118), .B1(new_n787), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n446), .B(new_n1120), .C1(G132), .C2(new_n793), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n784), .A2(new_n857), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G128), .A2(new_n796), .B1(new_n847), .B2(G50), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n812), .A2(G159), .B1(new_n775), .B2(G137), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n771), .B1(new_n1117), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1079), .B(new_n1128), .C1(new_n431), .C2(new_n843), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT116), .Z(new_n1130));
  AND2_X1   g0930(.A1(new_n1112), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n834), .C1(new_n703), .C2(new_n721), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n905), .B2(new_n912), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n951), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n935), .A2(new_n1134), .A3(new_n938), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n742), .A2(new_n686), .A3(new_n834), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n953), .B1(new_n905), .B2(new_n912), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n954), .A2(new_n913), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n1134), .B1(new_n949), .B2(new_n950), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1133), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1134), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1111), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1136), .A2(new_n953), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n913), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n1134), .A3(new_n935), .A4(new_n938), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1132), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n913), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1141), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1131), .B1(new_n1150), .B2(new_n749), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n916), .A2(new_n917), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n534), .A2(G330), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n946), .A2(new_n496), .A3(new_n651), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1147), .A2(new_n913), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n954), .B1(new_n1155), .B2(new_n1133), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n905), .A2(new_n912), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1132), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(new_n1148), .A3(new_n953), .A4(new_n1136), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1154), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT114), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(new_n1150), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1141), .A3(new_n1149), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n697), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1151), .B1(new_n1162), .B2(new_n1164), .ZN(G378));
  AND3_X1   g0965(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n935), .A2(new_n938), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n1167), .B2(new_n940), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n925), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n723), .B1(new_n939), .B2(new_n941), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n913), .A2(new_n918), .A3(new_n923), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n923), .B1(new_n913), .B2(new_n918), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n903), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1170), .B(new_n958), .C1(new_n1173), .C2(new_n881), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n644), .A2(new_n496), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n680), .B1(new_n483), .B2(new_n485), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1169), .A2(new_n1174), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1154), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1163), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1163), .B2(new_n1185), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1181), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n925), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n881), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n955), .B1(new_n922), .B2(new_n923), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1171), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n958), .B1(new_n1194), .B2(new_n1170), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1190), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1169), .A2(new_n1174), .A3(new_n1181), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1189), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n697), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1187), .A2(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n805), .A2(new_n258), .B1(new_n799), .B2(new_n429), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G97), .B2(new_n775), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n446), .A2(new_n374), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n788), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n850), .A2(new_n502), .B1(G107), .B2(new_n793), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n812), .A2(G68), .B1(new_n809), .B2(G77), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G50), .B1(new_n278), .B2(new_n374), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1207), .A2(new_n1208), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT117), .B(G124), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n788), .C2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(G159), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n850), .A2(G137), .B1(G128), .B2(new_n793), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n784), .B2(new_n1118), .ZN(new_n1215));
  INV_X1    g1015(.A(G132), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1119), .A2(new_n805), .B1(new_n803), .B2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G150), .C2(new_n812), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT59), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1212), .B1(new_n1213), .B2(new_n799), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1218), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1210), .B1(new_n1208), .B2(new_n1207), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1223), .A2(new_n764), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n750), .B1(new_n844), .B2(G50), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1190), .C2(new_n765), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1184), .B2(new_n749), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1200), .A2(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1157), .A2(new_n765), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n750), .B1(new_n844), .B2(G68), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n781), .A2(new_n202), .B1(new_n791), .B2(new_n857), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT123), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n446), .B1(new_n788), .B2(G128), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n858), .B2(new_n794), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n805), .A2(new_n1216), .B1(new_n799), .B2(new_n429), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n803), .A2(new_n1118), .B1(new_n784), .B2(new_n1213), .ZN(new_n1237));
  OR4_X1    g1037(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n796), .A2(G294), .B1(new_n850), .B2(G107), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n258), .B2(new_n803), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT121), .Z(new_n1241));
  AOI22_X1  g1041(.A1(new_n812), .A2(new_n502), .B1(G283), .B2(new_n793), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT122), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT122), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n446), .B1(new_n787), .B2(new_n782), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n981), .B(new_n1246), .C1(G97), .C2(new_n809), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1238), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1231), .B1(new_n1249), .B2(new_n764), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1229), .A2(new_n749), .B1(new_n1230), .B2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1031), .B(KEYINPUT120), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1229), .B2(new_n1185), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1161), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1151), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1161), .A2(new_n1150), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1164), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1073), .A2(new_n825), .A3(new_n1074), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1257), .A2(new_n1261), .A3(new_n1255), .A4(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n681), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1261), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  NOR2_X1   g1068(.A1(new_n1229), .A2(new_n1185), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1229), .A2(new_n1185), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(KEYINPUT60), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1156), .A2(new_n1159), .A3(new_n1154), .A4(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n697), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1251), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n842), .A3(new_n869), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G384), .B(new_n1251), .C1(new_n1271), .C2(new_n1273), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1266), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1196), .A2(new_n1282), .A3(new_n1197), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1281), .A2(new_n1283), .A3(new_n749), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1196), .A2(new_n1186), .A3(new_n1197), .A4(new_n1252), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1226), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1261), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1227), .C1(new_n1187), .C2(new_n1199), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1266), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1280), .B1(new_n1290), .B2(KEYINPUT126), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1287), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1281), .A2(new_n1283), .A3(new_n749), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1265), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n998), .B(G390), .C1(new_n1018), .C2(new_n1033), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1262), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1303), .A2(new_n1262), .A3(new_n1306), .A4(new_n1304), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1265), .B(new_n1300), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1299), .A2(new_n1301), .A3(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1310), .B1(new_n1290), .B2(new_n1280), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(KEYINPUT127), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1320), .B2(new_n1322), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1261), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1289), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1300), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1300), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1324), .A2(new_n1289), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1321), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1326), .A2(new_n1309), .A3(new_n1308), .A4(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(G402));
endmodule


