

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U551 ( .A1(KEYINPUT33), .A2(n756), .ZN(n787) );
  NOR2_X1 U552 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U553 ( .A(KEYINPUT29), .B(n717), .Z(n518) );
  AND2_X1 U554 ( .A1(n537), .A2(n536), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n798), .A2(n757), .ZN(n520) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n727) );
  XNOR2_X1 U557 ( .A(n727), .B(KEYINPUT102), .ZN(n728) );
  XNOR2_X1 U558 ( .A(n729), .B(n728), .ZN(n730) );
  INV_X1 U559 ( .A(n962), .ZN(n752) );
  NAND2_X1 U560 ( .A1(n692), .A2(n759), .ZN(n732) );
  AND2_X1 U561 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U562 ( .A1(n640), .A2(n526), .ZN(n646) );
  AND2_X2 U563 ( .A1(n538), .A2(G2104), .ZN(n893) );
  NOR2_X1 U564 ( .A1(n640), .A2(G651), .ZN(n655) );
  NOR2_X1 U565 ( .A1(G543), .A2(G651), .ZN(n649) );
  NAND2_X1 U566 ( .A1(G89), .A2(n649), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n521), .B(KEYINPUT74), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n522), .B(KEYINPUT4), .ZN(n524) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  INV_X1 U570 ( .A(G651), .ZN(n526) );
  NAND2_X1 U571 ( .A1(G76), .A2(n646), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n525), .B(KEYINPUT5), .ZN(n533) );
  NAND2_X1 U574 ( .A1(n655), .A2(G51), .ZN(n530) );
  NOR2_X1 U575 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n527), .Z(n528) );
  XNOR2_X1 U577 ( .A(KEYINPUT66), .B(n528), .ZN(n650) );
  NAND2_X1 U578 ( .A1(G63), .A2(n650), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n531), .Z(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U582 ( .A(n534), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  XOR2_X1 U585 ( .A(KEYINPUT17), .B(n535), .Z(n607) );
  NAND2_X1 U586 ( .A1(n607), .A2(G138), .ZN(n541) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U588 ( .A1(G114), .A2(n896), .ZN(n537) );
  NOR2_X1 U589 ( .A1(G2104), .A2(n538), .ZN(n605) );
  NAND2_X1 U590 ( .A1(G126), .A2(n605), .ZN(n536) );
  INV_X1 U591 ( .A(G2105), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G102), .A2(n893), .ZN(n539) );
  AND2_X1 U593 ( .A1(n519), .A2(n539), .ZN(n540) );
  AND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U595 ( .A1(n607), .A2(G137), .ZN(n688) );
  NAND2_X1 U596 ( .A1(G101), .A2(n893), .ZN(n542) );
  XNOR2_X1 U597 ( .A(KEYINPUT23), .B(n542), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G113), .A2(n896), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G125), .A2(n605), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n686) );
  AND2_X1 U602 ( .A1(n688), .A2(n686), .ZN(G160) );
  XOR2_X1 U603 ( .A(G2430), .B(G2451), .Z(n548) );
  XNOR2_X1 U604 ( .A(KEYINPUT109), .B(G2443), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n548), .B(n547), .ZN(n555) );
  XOR2_X1 U606 ( .A(G2435), .B(G2446), .Z(n550) );
  XNOR2_X1 U607 ( .A(G2427), .B(G2454), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(n551), .B(G2438), .Z(n553) );
  XNOR2_X1 U610 ( .A(G1341), .B(G1348), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n555), .B(n554), .ZN(n556) );
  AND2_X1 U613 ( .A1(n556), .A2(G14), .ZN(G401) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U619 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n834) );
  NAND2_X1 U621 ( .A1(n834), .A2(G567), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  NAND2_X1 U623 ( .A1(n650), .A2(G56), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n559), .Z(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT12), .B(KEYINPUT70), .Z(n561) );
  NAND2_X1 U626 ( .A1(G81), .A2(n649), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n646), .A2(G68), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT71), .B(n562), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT13), .ZN(n566) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n655), .A2(G43), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n973) );
  INV_X1 U635 ( .A(G860), .ZN(n623) );
  OR2_X1 U636 ( .A1(n973), .A2(n623), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G52), .A2(n655), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT68), .B(n570), .Z(n575) );
  NAND2_X1 U639 ( .A1(G90), .A2(n649), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G77), .A2(n646), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G64), .A2(n650), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U647 ( .A1(G92), .A2(n649), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n655), .A2(G54), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G66), .A2(n650), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n646), .A2(G79), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT72), .B(n580), .Z(n581) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT15), .ZN(n586) );
  XNOR2_X2 U655 ( .A(KEYINPUT73), .B(n586), .ZN(n978) );
  INV_X1 U656 ( .A(G868), .ZN(n668) );
  NAND2_X1 U657 ( .A1(n978), .A2(n668), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U659 ( .A1(n655), .A2(G53), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G65), .A2(n650), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G91), .A2(n649), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G78), .A2(n646), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n972) );
  XNOR2_X1 U666 ( .A(n972), .B(KEYINPUT69), .ZN(G299) );
  XNOR2_X1 U667 ( .A(KEYINPUT75), .B(G868), .ZN(n595) );
  NOR2_X1 U668 ( .A1(G286), .A2(n595), .ZN(n597) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n623), .A2(G559), .ZN(n598) );
  INV_X1 U672 ( .A(n978), .ZN(n621) );
  NAND2_X1 U673 ( .A1(n598), .A2(n621), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n973), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G868), .A2(n621), .ZN(n600) );
  NOR2_X1 U677 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G99), .A2(n893), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G111), .A2(n896), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n612) );
  BUF_X1 U682 ( .A(n605), .Z(n897) );
  NAND2_X1 U683 ( .A1(G123), .A2(n897), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT18), .ZN(n610) );
  BUF_X1 U685 ( .A(n607), .Z(n892) );
  NAND2_X1 U686 ( .A1(G135), .A2(n892), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT76), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n929) );
  XNOR2_X1 U690 ( .A(n929), .B(G2096), .ZN(n614) );
  INV_X1 U691 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n649), .A2(G93), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G67), .A2(n650), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G55), .A2(n655), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G80), .A2(n646), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n667) );
  NAND2_X1 U700 ( .A1(G559), .A2(n621), .ZN(n622) );
  XOR2_X1 U701 ( .A(n973), .B(n622), .Z(n665) );
  NAND2_X1 U702 ( .A1(n623), .A2(n665), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT77), .ZN(n625) );
  XOR2_X1 U704 ( .A(n667), .B(n625), .Z(G145) );
  NAND2_X1 U705 ( .A1(n655), .A2(G47), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G60), .A2(n650), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U708 ( .A(KEYINPUT67), .B(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G85), .A2(n649), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G72), .A2(n646), .ZN(n629) );
  AND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U713 ( .A1(n649), .A2(G88), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G62), .A2(n650), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G50), .A2(n655), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G75), .A2(n646), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n639), .Z(G166) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G87), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n650), .A2(n643), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n655), .A2(G49), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(G288) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n648) );
  NAND2_X1 U728 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n649), .A2(G86), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n655), .A2(G48), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(G305) );
  XNOR2_X1 U736 ( .A(G290), .B(G299), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U738 ( .A(G288), .B(KEYINPUT81), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(G166), .B(n660), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n667), .B(G305), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(n841) );
  XNOR2_X1 U744 ( .A(n841), .B(n665), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XOR2_X1 U749 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n671) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U757 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G96), .A2(n678), .ZN(n838) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n838), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT83), .B(n679), .ZN(n684) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G108), .A2(n681), .ZN(n839) );
  NAND2_X1 U764 ( .A1(G567), .A2(n839), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT84), .B(n682), .Z(n683) );
  NOR2_X1 U766 ( .A1(n684), .A2(n683), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n910) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n910), .A2(n685), .ZN(n837) );
  NAND2_X1 U770 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U771 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  INV_X1 U772 ( .A(G301), .ZN(G171) );
  AND2_X1 U773 ( .A1(n686), .A2(G40), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT87), .B(n689), .Z(n760) );
  INV_X1 U776 ( .A(n760), .ZN(n692) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n691) );
  INV_X1 U778 ( .A(KEYINPUT65), .ZN(n690) );
  XNOR2_X1 U779 ( .A(n691), .B(n690), .ZN(n759) );
  INV_X1 U780 ( .A(n732), .ZN(n704) );
  XOR2_X1 U781 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NAND2_X1 U782 ( .A1(n704), .A2(n948), .ZN(n694) );
  NAND2_X1 U783 ( .A1(G1961), .A2(n732), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U785 ( .A(KEYINPUT100), .B(n695), .Z(n719) );
  NAND2_X1 U786 ( .A1(n719), .A2(G171), .ZN(n718) );
  NAND2_X1 U787 ( .A1(n704), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U788 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U789 ( .A(G1956), .ZN(n992) );
  NOR2_X1 U790 ( .A1(n992), .A2(n704), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n712) );
  NOR2_X1 U792 ( .A1(n972), .A2(n712), .ZN(n699) );
  XOR2_X1 U793 ( .A(n699), .B(KEYINPUT28), .Z(n716) );
  AND2_X1 U794 ( .A1(n704), .A2(G1996), .ZN(n700) );
  XOR2_X1 U795 ( .A(n700), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U796 ( .A1(n732), .A2(G1341), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n973), .A2(n703), .ZN(n708) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n732), .ZN(n706) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n704), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n978), .A2(n709), .ZN(n707) );
  OR2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n978), .A2(n709), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n972), .A2(n712), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n518), .ZN(n731) );
  NOR2_X1 U810 ( .A1(G171), .A2(n719), .ZN(n726) );
  INV_X1 U811 ( .A(KEYINPUT101), .ZN(n721) );
  NAND2_X1 U812 ( .A1(G8), .A2(n732), .ZN(n798) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n798), .ZN(n743) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n732), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n720) );
  XNOR2_X1 U816 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U817 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U818 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U819 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n744) );
  NAND2_X1 U822 ( .A1(n744), .A2(G286), .ZN(n738) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n732), .ZN(n733) );
  XNOR2_X1 U824 ( .A(n733), .B(KEYINPUT104), .ZN(n735) );
  NOR2_X1 U825 ( .A1(n798), .A2(G1971), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U829 ( .A(KEYINPUT105), .B(n739), .Z(n740) );
  NAND2_X1 U830 ( .A1(G8), .A2(n740), .ZN(n741) );
  XNOR2_X1 U831 ( .A(n741), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U832 ( .A1(G8), .A2(n742), .ZN(n747) );
  XNOR2_X1 U833 ( .A(KEYINPUT103), .B(n744), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n743), .A2(n745), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n790) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n961) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NOR2_X1 U839 ( .A1(n961), .A2(n968), .ZN(n750) );
  XNOR2_X1 U840 ( .A(n750), .B(KEYINPUT106), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n790), .A2(n751), .ZN(n754) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NOR2_X1 U843 ( .A1(n798), .A2(n752), .ZN(n753) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT64), .ZN(n756) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n982) );
  INV_X1 U846 ( .A(n982), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n961), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n520), .ZN(n785) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT88), .ZN(n829) );
  INV_X1 U851 ( .A(n829), .ZN(n784) );
  NAND2_X1 U852 ( .A1(G131), .A2(n892), .ZN(n763) );
  NAND2_X1 U853 ( .A1(G107), .A2(n896), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G95), .A2(n893), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G119), .A2(n897), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  OR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n876) );
  NAND2_X1 U859 ( .A1(G1991), .A2(n876), .ZN(n768) );
  XNOR2_X1 U860 ( .A(n768), .B(KEYINPUT92), .ZN(n782) );
  XOR2_X1 U861 ( .A(KEYINPUT38), .B(KEYINPUT97), .Z(n770) );
  NAND2_X1 U862 ( .A1(G105), .A2(n893), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U864 ( .A(KEYINPUT96), .B(n771), .Z(n778) );
  NAND2_X1 U865 ( .A1(n897), .A2(G129), .ZN(n772) );
  XNOR2_X1 U866 ( .A(KEYINPUT93), .B(n772), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n896), .A2(G117), .ZN(n773) );
  XOR2_X1 U868 ( .A(KEYINPUT94), .B(n773), .Z(n774) );
  NOR2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U870 ( .A(KEYINPUT95), .B(n776), .ZN(n777) );
  NOR2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n892), .A2(G141), .ZN(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n874) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n874), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U876 ( .A(KEYINPUT98), .B(n783), .Z(n930) );
  NOR2_X1 U877 ( .A1(n784), .A2(n930), .ZN(n823) );
  INV_X1 U878 ( .A(n823), .ZN(n792) );
  AND2_X1 U879 ( .A1(n785), .A2(n792), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n803) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n788) );
  NAND2_X1 U882 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U884 ( .A(KEYINPUT107), .B(n791), .Z(n794) );
  AND2_X1 U885 ( .A1(n798), .A2(n792), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n801) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT99), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT24), .ZN(n797) );
  OR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U891 ( .A1(n823), .A2(n799), .ZN(n800) );
  AND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n819) );
  XOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .Z(n804) );
  XNOR2_X1 U895 ( .A(KEYINPUT89), .B(n804), .ZN(n827) );
  NAND2_X1 U896 ( .A1(G140), .A2(n892), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G104), .A2(n893), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n807), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G116), .A2(n896), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G128), .A2(n897), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT90), .B(n811), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(n814), .ZN(n906) );
  NOR2_X1 U907 ( .A1(n827), .A2(n906), .ZN(n815) );
  XNOR2_X1 U908 ( .A(n815), .B(KEYINPUT91), .ZN(n934) );
  XOR2_X1 U909 ( .A(G1986), .B(KEYINPUT86), .Z(n816) );
  XNOR2_X1 U910 ( .A(G290), .B(n816), .ZN(n971) );
  NAND2_X1 U911 ( .A1(n934), .A2(n971), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n829), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n832) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n874), .ZN(n922) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n876), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT108), .B(n820), .ZN(n933) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n933), .A2(n821), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n922), .A2(n824), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n934), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n906), .A2(n827), .ZN(n926) );
  NAND2_X1 U924 ( .A1(n828), .A2(n926), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(G286), .B(n973), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U942 ( .A(n978), .B(G171), .Z(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  NOR2_X1 U944 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U945 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U946 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U954 ( .A(KEYINPUT112), .B(G1976), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1956), .B(G1981), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U960 ( .A(G1971), .B(G1961), .Z(n860) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1966), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U964 ( .A(KEYINPUT111), .B(G2474), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n897), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G112), .A2(n896), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(n866), .Z(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G136), .A2(n892), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G100), .A2(n893), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U975 ( .A(G160), .B(n929), .Z(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U977 ( .A(G164), .B(G162), .Z(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(n878), .B(n877), .Z(n883) );
  XOR2_X1 U980 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT46), .B(n881), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n908) );
  NAND2_X1 U985 ( .A1(G142), .A2(n892), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G106), .A2(n893), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n886), .B(KEYINPUT45), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G118), .A2(n896), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G130), .A2(n897), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U992 ( .A(KEYINPUT114), .B(n889), .Z(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n904) );
  NAND2_X1 U994 ( .A1(G139), .A2(n892), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G115), .A2(n896), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(KEYINPUT117), .B(n903), .Z(n917) );
  XNOR2_X1 U1003 ( .A(n904), .B(n917), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n910), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n915), .A2(G395), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(KEYINPUT119), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1016 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n920), .Z(n925) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n938) );
  XOR2_X1 U1025 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n1016), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1036 ( .A(G2084), .B(G34), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(KEYINPUT54), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n958) );
  XOR2_X1 U1040 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n956) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1051 ( .A(n956), .B(n955), .Z(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n1017) );
  NOR2_X1 U1053 ( .A1(G29), .A2(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n1017), .A2(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n960), .ZN(n1023) );
  XOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .Z(n990) );
  INV_X1 U1057 ( .A(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT123), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(G1971), .A2(G303), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT124), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n988) );
  XNOR2_X1 U1065 ( .A(n972), .B(G1956), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G301), .B(G1961), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n973), .B(G1341), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1348), .B(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT122), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT57), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n991), .ZN(n1021) );
  XOR2_X1 U1080 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n1014) );
  XNOR2_X1 U1081 ( .A(G20), .B(n992), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1087 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(KEYINPUT60), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G1961), .B(G5), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1012) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT126), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(G16), .A2(n1015), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

