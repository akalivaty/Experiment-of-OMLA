

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U552 ( .A(n887), .Z(n516) );
  XOR2_X1 U553 ( .A(KEYINPUT17), .B(n536), .Z(n887) );
  XNOR2_X1 U554 ( .A(n653), .B(KEYINPUT91), .ZN(n640) );
  NOR2_X1 U555 ( .A1(G299), .A2(n634), .ZN(n602) );
  NOR2_X1 U556 ( .A1(n680), .A2(KEYINPUT33), .ZN(n682) );
  INV_X1 U557 ( .A(KEYINPUT97), .ZN(n681) );
  INV_X1 U558 ( .A(KEYINPUT92), .ZN(n601) );
  AND2_X1 U559 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U560 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U561 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NOR2_X1 U563 ( .A1(G651), .A2(n555), .ZN(n778) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n517) );
  XNOR2_X1 U565 ( .A(KEYINPUT64), .B(n517), .ZN(n555) );
  NAND2_X1 U566 ( .A1(n778), .A2(G53), .ZN(n519) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(G651), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n555), .A2(n520), .ZN(n774) );
  NAND2_X1 U569 ( .A1(G78), .A2(n774), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n773) );
  NAND2_X1 U572 ( .A1(n773), .A2(G91), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n522) );
  NOR2_X1 U574 ( .A1(G543), .A2(n520), .ZN(n521) );
  XNOR2_X1 U575 ( .A(n522), .B(n521), .ZN(n779) );
  NAND2_X1 U576 ( .A1(G65), .A2(n779), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n525) );
  OR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(G299) );
  NAND2_X1 U579 ( .A1(G86), .A2(n773), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G48), .A2(n778), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n774), .A2(G73), .ZN(n529) );
  XOR2_X1 U583 ( .A(KEYINPUT2), .B(n529), .Z(n530) );
  NOR2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G61), .A2(n779), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(G305) );
  INV_X1 U587 ( .A(G2105), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n537), .ZN(n878) );
  NAND2_X1 U589 ( .A1(G126), .A2(n878), .ZN(n535) );
  AND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U591 ( .A1(G114), .A2(n880), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n544) );
  NAND2_X1 U593 ( .A1(G138), .A2(n516), .ZN(n540) );
  AND2_X1 U594 ( .A1(n537), .A2(G2104), .ZN(n884) );
  NAND2_X1 U595 ( .A1(n884), .A2(G102), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT86), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n542) );
  INV_X1 U598 ( .A(KEYINPUT87), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n542), .B(n541), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n544), .A2(n543), .ZN(G164) );
  NAND2_X1 U601 ( .A1(n516), .A2(G137), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G101), .A2(n884), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(n545), .Z(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G125), .A2(n878), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G113), .A2(n880), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G160) );
  NAND2_X1 U609 ( .A1(G49), .A2(n778), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G74), .A2(G651), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n779), .A2(n554), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n555), .A2(G87), .ZN(n556) );
  XOR2_X1 U614 ( .A(KEYINPUT79), .B(n556), .Z(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(G288) );
  NAND2_X1 U616 ( .A1(n778), .A2(G52), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G64), .A2(n779), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U619 ( .A(KEYINPUT68), .B(n561), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n773), .A2(G90), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G77), .A2(n774), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(G171) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT72), .ZN(n578) );
  NAND2_X1 U626 ( .A1(n773), .A2(G89), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G76), .A2(n774), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U630 ( .A(KEYINPUT5), .B(n570), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G63), .A2(n779), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT71), .B(n571), .Z(n573) );
  NAND2_X1 U633 ( .A1(n778), .A2(G51), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U637 ( .A(n578), .B(n577), .ZN(G168) );
  NAND2_X1 U638 ( .A1(n778), .A2(G50), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G75), .A2(n774), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n773), .A2(G88), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT80), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G62), .A2(n779), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(G303) );
  INV_X1 U646 ( .A(G303), .ZN(G166) );
  XOR2_X1 U647 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U648 ( .A1(n773), .A2(G85), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G72), .A2(n774), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U651 ( .A(KEYINPUT66), .B(n588), .Z(n592) );
  NAND2_X1 U652 ( .A1(n779), .A2(G60), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n778), .A2(G47), .ZN(n589) );
  AND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(G290) );
  XOR2_X1 U656 ( .A(G1981), .B(G305), .Z(n961) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n699) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n698) );
  INV_X1 U659 ( .A(n698), .ZN(n593) );
  NAND2_X2 U660 ( .A1(n699), .A2(n593), .ZN(n653) );
  NAND2_X1 U661 ( .A1(G8), .A2(n653), .ZN(n693) );
  NOR2_X1 U662 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NAND2_X1 U663 ( .A1(n969), .A2(KEYINPUT33), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n693), .A2(n594), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT98), .B(n595), .Z(n596) );
  NAND2_X1 U666 ( .A1(n961), .A2(n596), .ZN(n684) );
  NAND2_X1 U667 ( .A1(n640), .A2(G2072), .ZN(n597) );
  XOR2_X1 U668 ( .A(KEYINPUT27), .B(n597), .Z(n600) );
  INV_X1 U669 ( .A(n640), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G1956), .A2(n598), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n634) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n633) );
  NAND2_X1 U673 ( .A1(G79), .A2(n774), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT70), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G54), .A2(n778), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n773), .A2(G92), .ZN(n607) );
  NAND2_X1 U678 ( .A1(G66), .A2(n779), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT69), .B(n608), .Z(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT15), .B(n611), .Z(n898) );
  NAND2_X1 U683 ( .A1(n779), .A2(G56), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT14), .B(n612), .Z(n618) );
  NAND2_X1 U685 ( .A1(n773), .A2(G81), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT12), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G68), .A2(n774), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U689 ( .A(KEYINPUT13), .B(n616), .Z(n617) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n778), .A2(G43), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n964) );
  INV_X1 U693 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U694 ( .A1(n653), .A2(n942), .ZN(n621) );
  XOR2_X1 U695 ( .A(n621), .B(KEYINPUT26), .Z(n623) );
  NAND2_X1 U696 ( .A1(n653), .A2(G1341), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n964), .A2(n624), .ZN(n625) );
  OR2_X1 U699 ( .A1(n898), .A2(n625), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n898), .A2(n625), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G2067), .A2(n640), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G1348), .A2(n653), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U707 ( .A1(G299), .A2(n634), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT28), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U710 ( .A(KEYINPUT93), .B(KEYINPUT29), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n644) );
  INV_X1 U712 ( .A(G1961), .ZN(n913) );
  NAND2_X1 U713 ( .A1(n913), .A2(n653), .ZN(n642) );
  XNOR2_X1 U714 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NAND2_X1 U715 ( .A1(n640), .A2(n941), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n649), .A2(G171), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n667) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n693), .ZN(n669) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n653), .ZN(n665) );
  NOR2_X1 U721 ( .A1(n669), .A2(n665), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G8), .A2(n645), .ZN(n647) );
  XNOR2_X1 U723 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U725 ( .A1(G168), .A2(n648), .ZN(n651) );
  NOR2_X1 U726 ( .A1(G171), .A2(n649), .ZN(n650) );
  NOR2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U728 ( .A(KEYINPUT31), .B(n652), .Z(n666) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(KEYINPUT95), .B(n654), .ZN(n657) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n693), .ZN(n655) );
  NOR2_X1 U732 ( .A1(G166), .A2(n655), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n659) );
  AND2_X1 U734 ( .A1(n666), .A2(n659), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n667), .A2(n658), .ZN(n662) );
  INV_X1 U736 ( .A(n659), .ZN(n660) );
  OR2_X1 U737 ( .A1(n660), .A2(G286), .ZN(n661) );
  AND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n663), .A2(G8), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(KEYINPUT32), .ZN(n673) );
  NAND2_X1 U741 ( .A1(G8), .A2(n665), .ZN(n671) );
  AND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U743 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n686) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n674) );
  NOR2_X1 U747 ( .A1(n969), .A2(n674), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n686), .A2(n675), .ZN(n679) );
  INV_X1 U749 ( .A(n693), .ZN(n677) );
  NAND2_X1 U750 ( .A1(G288), .A2(G1976), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n676), .B(KEYINPUT96), .ZN(n970) );
  AND2_X1 U752 ( .A1(n677), .A2(n970), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT99), .ZN(n697) );
  NOR2_X1 U754 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U755 ( .A1(G8), .A2(n687), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n686), .A2(n688), .ZN(n689) );
  AND2_X1 U757 ( .A1(n689), .A2(n693), .ZN(n695) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U759 ( .A(n690), .B(KEYINPUT90), .Z(n691) );
  XNOR2_X1 U760 ( .A(KEYINPUT24), .B(n691), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n731) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n743) );
  XNOR2_X1 U765 ( .A(KEYINPUT37), .B(G2067), .ZN(n732) );
  NAND2_X1 U766 ( .A1(n516), .A2(G140), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U768 ( .A1(G104), .A2(n884), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(KEYINPUT34), .B(n703), .ZN(n708) );
  NAND2_X1 U771 ( .A1(G128), .A2(n878), .ZN(n705) );
  NAND2_X1 U772 ( .A1(G116), .A2(n880), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U774 ( .A(KEYINPUT35), .B(n706), .Z(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(KEYINPUT36), .B(n709), .ZN(n895) );
  NOR2_X1 U777 ( .A1(n732), .A2(n895), .ZN(n1009) );
  NAND2_X1 U778 ( .A1(n743), .A2(n1009), .ZN(n739) );
  NAND2_X1 U779 ( .A1(G95), .A2(n884), .ZN(n711) );
  NAND2_X1 U780 ( .A1(G131), .A2(n516), .ZN(n710) );
  NAND2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G119), .A2(n878), .ZN(n713) );
  NAND2_X1 U783 ( .A1(G107), .A2(n880), .ZN(n712) );
  NAND2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n861) );
  INV_X1 U786 ( .A(G1991), .ZN(n937) );
  NOR2_X1 U787 ( .A1(n861), .A2(n937), .ZN(n725) );
  NAND2_X1 U788 ( .A1(G141), .A2(n516), .ZN(n717) );
  NAND2_X1 U789 ( .A1(G129), .A2(n878), .ZN(n716) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U791 ( .A1(G105), .A2(n884), .ZN(n718) );
  XNOR2_X1 U792 ( .A(n718), .B(KEYINPUT38), .ZN(n719) );
  XNOR2_X1 U793 ( .A(n719), .B(KEYINPUT89), .ZN(n720) );
  NOR2_X1 U794 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n880), .A2(G117), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n892) );
  AND2_X1 U797 ( .A1(n892), .A2(G1996), .ZN(n724) );
  NOR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n994) );
  INV_X1 U799 ( .A(n743), .ZN(n726) );
  NOR2_X1 U800 ( .A1(n994), .A2(n726), .ZN(n735) );
  INV_X1 U801 ( .A(n735), .ZN(n727) );
  AND2_X1 U802 ( .A1(n739), .A2(n727), .ZN(n729) );
  XNOR2_X1 U803 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U804 ( .A1(n981), .A2(n743), .ZN(n728) );
  AND2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n746) );
  NAND2_X1 U807 ( .A1(n732), .A2(n895), .ZN(n1006) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n892), .ZN(n991) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n733) );
  AND2_X1 U810 ( .A1(n937), .A2(n861), .ZN(n989) );
  NOR2_X1 U811 ( .A1(n733), .A2(n989), .ZN(n734) );
  NOR2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U813 ( .A1(n991), .A2(n736), .ZN(n737) );
  XNOR2_X1 U814 ( .A(KEYINPUT100), .B(n737), .ZN(n738) );
  XNOR2_X1 U815 ( .A(n738), .B(KEYINPUT39), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n1006), .A2(n741), .ZN(n742) );
  XOR2_X1 U818 ( .A(KEYINPUT101), .B(n742), .Z(n744) );
  NAND2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U822 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U823 ( .A(G132), .ZN(G219) );
  INV_X1 U824 ( .A(G82), .ZN(G220) );
  INV_X1 U825 ( .A(G57), .ZN(G237) );
  NAND2_X1 U826 ( .A1(G7), .A2(G661), .ZN(n748) );
  XNOR2_X1 U827 ( .A(n748), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U828 ( .A(G223), .ZN(n825) );
  NAND2_X1 U829 ( .A1(n825), .A2(G567), .ZN(n749) );
  XOR2_X1 U830 ( .A(KEYINPUT11), .B(n749), .Z(G234) );
  INV_X1 U831 ( .A(G860), .ZN(n754) );
  OR2_X1 U832 ( .A1(n964), .A2(n754), .ZN(G153) );
  INV_X1 U833 ( .A(G171), .ZN(G301) );
  NAND2_X1 U834 ( .A1(G868), .A2(G301), .ZN(n751) );
  INV_X1 U835 ( .A(n898), .ZN(n975) );
  INV_X1 U836 ( .A(G868), .ZN(n757) );
  NAND2_X1 U837 ( .A1(n975), .A2(n757), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(G284) );
  NAND2_X1 U839 ( .A1(G868), .A2(G286), .ZN(n753) );
  NAND2_X1 U840 ( .A1(G299), .A2(n757), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(G297) );
  NAND2_X1 U842 ( .A1(n754), .A2(G559), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n755), .A2(n898), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U845 ( .A1(G559), .A2(n757), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n898), .A2(n758), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT73), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n964), .A2(G868), .ZN(n760) );
  NOR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(G282) );
  XOR2_X1 U850 ( .A(G2100), .B(KEYINPUT76), .Z(n772) );
  NAND2_X1 U851 ( .A1(G123), .A2(n878), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT74), .ZN(n763) );
  XNOR2_X1 U853 ( .A(KEYINPUT18), .B(n763), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G99), .A2(n884), .ZN(n764) );
  XOR2_X1 U855 ( .A(KEYINPUT75), .B(n764), .Z(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G135), .A2(n516), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G111), .A2(n880), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n988) );
  XNOR2_X1 U861 ( .A(G2096), .B(n988), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(G156) );
  NAND2_X1 U863 ( .A1(n773), .A2(G93), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G80), .A2(n774), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(KEYINPUT78), .B(n777), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n778), .A2(G55), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G67), .A2(n779), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n790) );
  NAND2_X1 U871 ( .A1(G559), .A2(n898), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(n964), .ZN(n794) );
  XOR2_X1 U873 ( .A(KEYINPUT77), .B(n794), .Z(n785) );
  NOR2_X1 U874 ( .A1(G860), .A2(n785), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n790), .B(n786), .ZN(G145) );
  NOR2_X1 U876 ( .A1(G868), .A2(n790), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(KEYINPUT81), .ZN(n797) );
  XNOR2_X1 U878 ( .A(KEYINPUT19), .B(G305), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(G288), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n790), .B(n789), .ZN(n792) );
  XNOR2_X1 U881 ( .A(G299), .B(G166), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n792), .B(n791), .ZN(n793) );
  XOR2_X1 U883 ( .A(n793), .B(G290), .Z(n899) );
  XNOR2_X1 U884 ( .A(n899), .B(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G868), .A2(n795), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(G295) );
  NAND2_X1 U887 ( .A1(G2078), .A2(G2084), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT20), .B(n798), .Z(n799) );
  NAND2_X1 U889 ( .A1(G2090), .A2(n799), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n801), .B(n800), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n802), .A2(G2072), .ZN(n803) );
  XOR2_X1 U893 ( .A(KEYINPUT83), .B(n803), .Z(G158) );
  XNOR2_X1 U894 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U895 ( .A1(G69), .A2(G120), .ZN(n804) );
  NOR2_X1 U896 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G108), .A2(n805), .ZN(n832) );
  NAND2_X1 U898 ( .A1(G567), .A2(n832), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT84), .ZN(n811) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n807) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n807), .Z(n808) );
  NOR2_X1 U902 ( .A1(G218), .A2(n808), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G96), .A2(n809), .ZN(n831) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n831), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U906 ( .A(KEYINPUT85), .B(n812), .ZN(G319) );
  INV_X1 U907 ( .A(G319), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G661), .A2(G483), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n830) );
  NAND2_X1 U910 ( .A1(n830), .A2(G36), .ZN(G176) );
  XNOR2_X1 U911 ( .A(G2430), .B(G2454), .ZN(n823) );
  XNOR2_X1 U912 ( .A(KEYINPUT102), .B(G2435), .ZN(n821) );
  XOR2_X1 U913 ( .A(G2451), .B(G2427), .Z(n816) );
  XNOR2_X1 U914 ( .A(G2438), .B(G2446), .ZN(n815) );
  XNOR2_X1 U915 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U916 ( .A(n817), .B(G2443), .Z(n819) );
  XNOR2_X1 U917 ( .A(G1341), .B(G1348), .ZN(n818) );
  XNOR2_X1 U918 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U919 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(G14), .ZN(n907) );
  XNOR2_X1 U922 ( .A(KEYINPUT103), .B(n907), .ZN(G401) );
  NAND2_X1 U923 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n826), .B(KEYINPUT104), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n827) );
  XNOR2_X1 U926 ( .A(KEYINPUT105), .B(n827), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n828), .A2(G661), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U929 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U930 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n833), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U936 ( .A(G261), .ZN(G325) );
  XOR2_X1 U937 ( .A(G2096), .B(G2100), .Z(n835) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n834) );
  XNOR2_X1 U939 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n837) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U942 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U943 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U945 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1966), .Z(n843) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U948 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U949 ( .A(n844), .B(KEYINPUT108), .Z(n846) );
  XNOR2_X1 U950 ( .A(G1956), .B(G1976), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U952 ( .A(G1981), .B(G1971), .Z(n848) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n847) );
  XNOR2_X1 U954 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U955 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(G2474), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G124), .A2(n878), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n853), .B(KEYINPUT44), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n854), .B(KEYINPUT110), .ZN(n856) );
  NAND2_X1 U961 ( .A1(G100), .A2(n884), .ZN(n855) );
  NAND2_X1 U962 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G136), .A2(n516), .ZN(n858) );
  NAND2_X1 U964 ( .A1(G112), .A2(n880), .ZN(n857) );
  NAND2_X1 U965 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U966 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n863) );
  XNOR2_X1 U968 ( .A(n861), .B(KEYINPUT112), .ZN(n862) );
  XNOR2_X1 U969 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U970 ( .A(n864), .B(n988), .Z(n866) );
  XNOR2_X1 U971 ( .A(G164), .B(G160), .ZN(n865) );
  XNOR2_X1 U972 ( .A(n866), .B(n865), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G106), .A2(n884), .ZN(n868) );
  NAND2_X1 U974 ( .A1(G142), .A2(n516), .ZN(n867) );
  NAND2_X1 U975 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U976 ( .A(n869), .B(KEYINPUT45), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G130), .A2(n878), .ZN(n871) );
  NAND2_X1 U978 ( .A1(G118), .A2(n880), .ZN(n870) );
  NAND2_X1 U979 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U980 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  NAND2_X1 U981 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U982 ( .A(n875), .B(G162), .ZN(n876) );
  XOR2_X1 U983 ( .A(n877), .B(n876), .Z(n894) );
  NAND2_X1 U984 ( .A1(n878), .A2(G127), .ZN(n879) );
  XNOR2_X1 U985 ( .A(n879), .B(KEYINPUT114), .ZN(n882) );
  NAND2_X1 U986 ( .A1(G115), .A2(n880), .ZN(n881) );
  NAND2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U988 ( .A(n883), .B(KEYINPUT47), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G103), .A2(n884), .ZN(n885) );
  NAND2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G139), .A2(n516), .ZN(n888) );
  XNOR2_X1 U992 ( .A(KEYINPUT113), .B(n888), .ZN(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(n891), .Z(n1000) );
  XOR2_X1 U995 ( .A(n892), .B(n1000), .Z(n893) );
  XNOR2_X1 U996 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U998 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U999 ( .A(KEYINPUT116), .B(n964), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n898), .B(G171), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(n903), .B(G286), .Z(n904) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n904), .ZN(G397) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n907), .ZN(n908) );
  XOR2_X1 U1009 ( .A(KEYINPUT117), .B(n908), .Z(n909) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(G5), .B(n913), .ZN(n930) );
  XOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .Z(n914) );
  XNOR2_X1 U1017 ( .A(G4), .B(n914), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(G20), .B(G1956), .ZN(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(G1981), .B(G6), .ZN(n917) );
  NOR2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(n921), .B(KEYINPUT60), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G1971), .B(G22), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(G23), .B(G1976), .ZN(n922) );
  NOR2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n925) );
  XOR2_X1 U1028 ( .A(G1986), .B(G24), .Z(n924) );
  NAND2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1030 ( .A(KEYINPUT58), .B(n926), .ZN(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G21), .B(G1966), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT61), .B(n933), .ZN(n935) );
  INV_X1 U1036 ( .A(G16), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n936), .A2(G11), .ZN(n1019) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n956) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(G25), .B(n937), .ZN(n938) );
  NAND2_X1 U1042 ( .A1(n938), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1045 ( .A1(n940), .A2(n939), .ZN(n946) );
  XOR2_X1 U1046 ( .A(n941), .B(G27), .Z(n944) );
  XOR2_X1 U1047 ( .A(n942), .B(G32), .Z(n943) );
  NOR2_X1 U1048 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n952) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n952), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n956), .B(n955), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(KEYINPUT55), .B(n957), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(G29), .B(KEYINPUT122), .ZN(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(KEYINPUT123), .B(n960), .ZN(n1017) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1063 ( .A(KEYINPUT57), .B(n963), .Z(n984) );
  XNOR2_X1 U1064 ( .A(n964), .B(G1341), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(G301), .B(G1961), .ZN(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G299), .B(G1956), .ZN(n968) );
  XNOR2_X1 U1068 ( .A(G303), .B(G1971), .ZN(n967) );
  NOR2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n974) );
  INV_X1 U1070 ( .A(n969), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1072 ( .A(KEYINPUT124), .B(n972), .Z(n973) );
  NAND2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n975), .ZN(n976) );
  NOR2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(KEYINPUT125), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .Z(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n987), .ZN(n1015) );
  INV_X1 U1083 ( .A(G29), .ZN(n1013) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n999) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(n992), .B(KEYINPUT119), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n993), .B(KEYINPUT51), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1090 ( .A(G160), .B(G2084), .Z(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1003), .Z(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1010), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(KEYINPUT55), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT127), .B(n1020), .Z(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

