//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G250), .B(G257), .Z(new_n225));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  AND2_X1   g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NOR2_X1   g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n247), .A2(G223), .B1(G77), .B2(new_n245), .ZN(new_n248));
  INV_X1    g0048(.A(G222), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n246), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n248), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n209), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G33), .A3(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(new_n257), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(G274), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(KEYINPUT68), .A2(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT68), .A2(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n265), .A2(new_n273), .A3(G226), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n261), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(G179), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT69), .B1(new_n203), .B2(new_n251), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n209), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n251), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n281), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G50), .A2(G58), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n210), .B1(new_n288), .B2(new_n214), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n280), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT68), .A2(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT68), .A2(G1), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n280), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n290), .B(new_n297), .C1(new_n296), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n275), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n276), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n275), .A2(G200), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n307), .B1(new_n306), .B2(new_n301), .C1(new_n308), .C2(new_n275), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n295), .A2(KEYINPUT12), .A3(new_n214), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT12), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n294), .B2(G68), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n283), .A2(new_n318), .B1(new_n210), .B2(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n286), .A2(new_n296), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n280), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n322), .B1(new_n317), .B2(new_n321), .C1(new_n214), .C2(new_n300), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  INV_X1    g0124(.A(G226), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n255), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n246), .A2(KEYINPUT72), .A3(G226), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n246), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n254), .B1(G33), .B2(G97), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n259), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n265), .A2(new_n273), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n269), .B1(new_n332), .B2(new_n215), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT13), .B1(new_n331), .B2(new_n333), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n338));
  OR3_X1    g0138(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n323), .B1(new_n340), .B2(G190), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(KEYINPUT73), .A3(new_n337), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT73), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n334), .A2(new_n343), .A3(new_n335), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(G200), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(G169), .A3(new_n344), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(G179), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n342), .A2(new_n350), .A3(G169), .A4(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n323), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G244), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n269), .B1(new_n332), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n245), .A2(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G232), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT70), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n247), .A2(G238), .B1(G107), .B2(new_n245), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n356), .B1(new_n361), .B2(new_n259), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n302), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n356), .C1(new_n361), .C2(new_n259), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G20), .A2(G77), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n281), .B2(new_n286), .C1(new_n283), .C2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n280), .B1(new_n295), .B2(new_n318), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n298), .A2(G77), .A3(new_n299), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n363), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n362), .A2(G200), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n370), .B(new_n369), .C1(new_n362), .C2(new_n308), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n312), .A2(new_n353), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n295), .A2(new_n281), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n300), .B2(new_n281), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n252), .A2(new_n210), .A3(new_n253), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n383), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n386), .B(G68), .C1(new_n389), .C2(new_n385), .ZN(new_n390));
  INV_X1    g0190(.A(G58), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n214), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n285), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT16), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n245), .B2(new_n210), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n384), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n280), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n381), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n265), .A2(new_n273), .A3(G232), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT76), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT76), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n265), .A2(new_n273), .A3(new_n407), .A4(G232), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n325), .A2(G1698), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G223), .B2(G1698), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n411), .A2(new_n245), .B1(new_n251), .B2(new_n216), .ZN(new_n412));
  INV_X1    g0212(.A(G274), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n209), .B1(KEYINPUT67), .B2(new_n258), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n264), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n412), .A2(new_n260), .B1(new_n415), .B2(new_n268), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(G190), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n325), .B2(G1698), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n254), .B1(G33), .B2(G87), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n269), .B1(new_n420), .B2(new_n259), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n408), .B2(new_n406), .ZN(new_n422));
  INV_X1    g0222(.A(G200), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n404), .A2(KEYINPUT17), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n403), .B2(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT77), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n409), .A2(new_n430), .A3(new_n416), .A4(new_n364), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n409), .A2(new_n364), .A3(new_n416), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n433));
  AOI21_X1  g0233(.A(G169), .B1(new_n409), .B2(new_n416), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT18), .B1(new_n435), .B2(new_n403), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n437), .A3(new_n436), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n429), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n378), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n299), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(G13), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT83), .B(KEYINPUT25), .C1(new_n294), .C2(G107), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n293), .A2(G33), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n298), .A2(new_n294), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(G107), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n210), .B(G87), .C1(new_n243), .C2(new_n244), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT22), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n254), .A2(new_n458), .A3(new_n210), .A4(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT23), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n210), .B2(G107), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n447), .A2(KEYINPUT23), .A3(G20), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n463), .A2(new_n464), .B1(new_n282), .B2(G116), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n460), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n461), .B1(new_n460), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n280), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n455), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n470));
  OAI211_X1 g0270(.A(G250), .B(new_n246), .C1(new_n243), .C2(new_n244), .ZN(new_n471));
  INV_X1    g0271(.A(G294), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n251), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n270), .A2(G45), .A3(new_n272), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n473), .A2(new_n260), .B1(new_n415), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n265), .B(G264), .C1(new_n474), .C2(new_n477), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n479), .B(G179), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n302), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI211_X1 g0286(.A(KEYINPUT84), .B(new_n302), .C1(new_n479), .C2(new_n480), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n469), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT86), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n480), .B(KEYINPUT85), .ZN(new_n491));
  AOI21_X1  g0291(.A(G200), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n479), .A2(new_n308), .A3(new_n480), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n468), .B(new_n455), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n469), .B(KEYINPUT86), .C1(new_n486), .C2(new_n487), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n490), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n245), .A2(G303), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n246), .C1(new_n243), .C2(new_n244), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G264), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n254), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n259), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n293), .B(G45), .C1(new_n476), .C2(new_n475), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G270), .A3(new_n265), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n478), .A2(new_n415), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(G169), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n298), .A2(G116), .A3(new_n294), .A4(new_n452), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n295), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(G33), .B2(G283), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n251), .A2(G97), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(G20), .B2(new_n514), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n280), .A2(KEYINPUT20), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT20), .B1(new_n280), .B2(new_n518), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n513), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n497), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n507), .A2(new_n511), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G179), .A3(new_n521), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n510), .B(new_n509), .C1(new_n526), .C2(new_n259), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(KEYINPUT21), .A3(G169), .A4(new_n521), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n523), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n521), .B1(new_n527), .B2(G200), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n308), .B2(new_n527), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n294), .A2(G97), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n453), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n386), .B(G107), .C1(new_n389), .C2(new_n385), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n447), .A2(KEYINPUT6), .A3(G97), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n536), .A2(new_n447), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(KEYINPUT6), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n533), .B(new_n538), .C1(new_n546), .C2(new_n298), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n254), .A2(G244), .A3(new_n246), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT4), .B1(new_n357), .B2(G244), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n260), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n508), .A2(G257), .A3(new_n265), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n555), .A2(new_n510), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n556), .A3(new_n308), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n510), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n357), .A2(KEYINPUT4), .A3(G244), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n548), .A4(new_n549), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n561), .B2(new_n260), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n557), .B1(new_n562), .B2(G200), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n298), .B1(new_n539), .B2(new_n545), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT79), .B1(new_n564), .B2(new_n537), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n547), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(G179), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n554), .A2(new_n556), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G169), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n538), .B1(new_n546), .B2(new_n298), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n254), .A2(G244), .A3(G1698), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n255), .C2(new_n215), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n260), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n270), .A2(G45), .A3(new_n413), .A4(new_n272), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n291), .A2(new_n292), .A3(new_n267), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n265), .B(new_n578), .C1(new_n579), .C2(G250), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G190), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n423), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n210), .B(G68), .C1(new_n243), .C2(new_n244), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n216), .A2(new_n536), .A3(new_n447), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT80), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G87), .A2(G97), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n447), .ZN(new_n596));
  NAND3_X1  g0396(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n593), .A2(new_n596), .B1(new_n210), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n280), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n367), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n294), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n298), .A2(G87), .A3(new_n294), .A4(new_n452), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n210), .ZN(new_n605));
  NOR4_X1   g0405(.A1(KEYINPUT80), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n595), .B1(new_n594), .B2(new_n447), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(new_n589), .A3(new_n590), .A4(new_n587), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n601), .B1(new_n609), .B2(new_n280), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n367), .B2(new_n453), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n577), .A2(new_n580), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(G179), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n581), .A2(G169), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n583), .A2(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n532), .A2(new_n573), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n445), .A2(new_n496), .A3(new_n616), .ZN(G372));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n580), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n474), .A2(new_n217), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(KEYINPUT87), .A3(new_n265), .A4(new_n578), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n622), .B2(new_n577), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n488), .A2(new_n523), .A3(new_n525), .A4(new_n528), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(new_n494), .A3(new_n572), .A4(new_n566), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n577), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT88), .B1(new_n610), .B2(new_n603), .ZN(new_n630));
  AND4_X1   g0430(.A1(KEYINPUT88), .A2(new_n599), .A3(new_n602), .A4(new_n603), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n627), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n582), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT88), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n604), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n610), .A2(KEYINPUT88), .A3(new_n603), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n627), .B1(new_n637), .B2(new_n629), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n624), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n624), .B1(new_n626), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n547), .A2(new_n565), .B1(new_n569), .B2(new_n567), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n624), .B(new_n641), .C1(new_n633), .C2(new_n638), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n615), .A2(new_n572), .ZN(new_n644));
  XNOR2_X1  g0444(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n642), .A2(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n445), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT92), .ZN(new_n650));
  INV_X1    g0450(.A(new_n429), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n341), .A2(new_n345), .ZN(new_n652));
  INV_X1    g0452(.A(new_n372), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n652), .A2(new_n653), .B1(new_n352), .B2(new_n323), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n352), .A2(new_n323), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(new_n658), .A3(new_n655), .ZN(new_n659));
  INV_X1    g0459(.A(new_n436), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n656), .A2(new_n659), .B1(new_n439), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n310), .A2(new_n311), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n650), .B1(new_n663), .B2(new_n304), .ZN(new_n664));
  AOI211_X1 g0464(.A(KEYINPUT92), .B(new_n305), .C1(new_n661), .C2(new_n662), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n649), .B1(new_n664), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n293), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G343), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n529), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n469), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n496), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n488), .B2(new_n674), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n488), .A2(new_n675), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  INV_X1    g0485(.A(new_n529), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n674), .A2(new_n522), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT93), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n532), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT95), .Z(G399));
  NOR2_X1   g0494(.A1(new_n606), .A2(new_n607), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n514), .ZN(new_n696));
  INV_X1    g0496(.A(G1), .ZN(new_n697));
  INV_X1    g0497(.A(new_n204), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n700), .A2(KEYINPUT96), .B1(new_n208), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(KEYINPUT96), .B2(new_n700), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n648), .A2(new_n674), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n645), .B1(new_n615), .B2(new_n572), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n642), .B2(new_n643), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n613), .A2(new_n623), .ZN(new_n709));
  INV_X1    g0509(.A(new_n582), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n635), .A2(new_n636), .B1(G200), .B2(new_n628), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n627), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n637), .A2(new_n629), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n566), .A2(new_n572), .A3(new_n494), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n490), .A2(new_n529), .A3(new_n495), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n708), .A2(new_n624), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n674), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n706), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n473), .A2(new_n260), .ZN(new_n723));
  AND4_X1   g0523(.A1(new_n723), .A2(new_n562), .A3(new_n581), .A4(new_n491), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n527), .A2(new_n364), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT98), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n724), .A2(new_n725), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n491), .A2(new_n479), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n568), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n527), .A2(new_n628), .A3(new_n364), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n729), .A2(KEYINPUT30), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n675), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n616), .A2(new_n496), .A3(new_n674), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT31), .B(new_n675), .C1(new_n728), .C2(new_n734), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n722), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n703), .B1(new_n742), .B2(new_n697), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT99), .Z(G364));
  AOI21_X1  g0544(.A(new_n209), .B1(G20), .B2(new_n302), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT100), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n698), .A2(new_n254), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n267), .B2(new_n208), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n238), .B2(new_n267), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n698), .A2(new_n245), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n514), .B2(new_n698), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n753), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n697), .B1(new_n668), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n699), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n210), .A2(new_n364), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n254), .B1(new_n767), .B2(new_n318), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n308), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n210), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n296), .B1(new_n216), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n766), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n768), .B(new_n774), .C1(KEYINPUT32), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n308), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n765), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT101), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G58), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n772), .A2(new_n308), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT102), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n447), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n777), .A2(KEYINPUT32), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n779), .A2(new_n364), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n536), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n769), .A2(G190), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n795), .B(new_n799), .C1(G68), .C2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n778), .A2(new_n787), .A3(new_n794), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G329), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n245), .B1(new_n775), .B2(new_n803), .C1(new_n804), .C2(new_n767), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n786), .B2(G322), .ZN(new_n806));
  INV_X1    g0606(.A(new_n792), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G283), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n770), .A2(G326), .B1(new_n797), .B2(G294), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  INV_X1    g0610(.A(new_n773), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n800), .A2(new_n810), .B1(new_n811), .B2(G303), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n806), .A2(new_n808), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n760), .B(new_n764), .C1(new_n814), .C2(new_n748), .ZN(new_n815));
  INV_X1    g0615(.A(new_n751), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n690), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n691), .A2(new_n764), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n690), .A2(G330), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT103), .Z(G396));
  AOI21_X1  g0621(.A(new_n245), .B1(new_n776), .B2(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n296), .B2(new_n773), .C1(new_n391), .C2(new_n798), .ZN(new_n823));
  INV_X1    g0623(.A(new_n767), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n770), .A2(G137), .B1(new_n824), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(new_n800), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n284), .B2(new_n826), .C1(new_n785), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  AOI211_X1 g0629(.A(new_n823), .B(new_n829), .C1(G68), .C2(new_n807), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n245), .B1(new_n775), .B2(new_n804), .C1(new_n514), .C2(new_n767), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n786), .B2(G294), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n799), .B1(G283), .B2(new_n800), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n770), .A2(G303), .B1(new_n811), .B2(G107), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G87), .B2(new_n807), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n748), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n748), .A2(new_n749), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n763), .C1(G77), .C2(new_n839), .ZN(new_n840));
  AND4_X1   g0640(.A1(new_n365), .A2(new_n363), .A3(new_n371), .A4(new_n674), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n675), .A2(new_n371), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n374), .B2(new_n373), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n372), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n840), .B1(new_n749), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n704), .A2(new_n845), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n674), .B(new_n844), .C1(new_n640), .C2(new_n647), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n763), .B1(new_n849), .B2(new_n741), .ZN(new_n850));
  INV_X1    g0650(.A(new_n741), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n847), .A3(new_n848), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  NOR2_X1   g0654(.A1(new_n293), .A2(new_n668), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n706), .A2(new_n445), .A3(new_n721), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n664), .B2(new_n665), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT109), .Z(new_n858));
  AOI21_X1  g0658(.A(new_n396), .B1(new_n389), .B2(G68), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n298), .B1(new_n859), .B2(KEYINPUT16), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT16), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n214), .B1(new_n387), .B2(new_n388), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n396), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n380), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n403), .A2(new_n424), .B1(new_n864), .B2(new_n672), .ZN(new_n865));
  OAI211_X1 g0665(.A(KEYINPUT77), .B(new_n432), .C1(new_n422), .C2(G169), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n866), .B2(new_n431), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n403), .B1(new_n435), .B2(new_n673), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n404), .A2(new_n425), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(KEYINPUT37), .C1(new_n865), .C2(new_n867), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n864), .A2(new_n672), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n443), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n876), .B(KEYINPUT38), .C1(new_n443), .C2(new_n877), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n841), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n848), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n323), .B(new_n675), .C1(new_n346), .C2(new_n352), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n323), .A2(new_n675), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n658), .A2(new_n652), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n882), .B1(new_n889), .B2(KEYINPUT104), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(KEYINPUT104), .B2(new_n889), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n660), .A2(new_n439), .A3(new_n673), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(new_n881), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n428), .B(new_n426), .C1(new_n660), .C2(new_n439), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n403), .A2(new_n673), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n872), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n435), .A2(new_n403), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n896), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n900), .B2(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n870), .A2(new_n871), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n895), .A2(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT108), .A4(new_n898), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n893), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT107), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n658), .B2(new_n675), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n352), .A2(KEYINPUT107), .A3(new_n323), .A4(new_n674), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n892), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n891), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n858), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n845), .B1(new_n885), .B2(new_n887), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n740), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n894), .A2(new_n905), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT40), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n882), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G330), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n851), .A2(new_n445), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT110), .Z(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n445), .A3(new_n740), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n855), .B1(new_n916), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n916), .B2(new_n928), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n211), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n392), .A2(new_n207), .A3(new_n318), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n296), .B2(G68), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n936), .A2(G13), .A3(new_n293), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  AOI21_X1  g0738(.A(new_n674), .B1(new_n547), .B2(new_n565), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n573), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n641), .A2(new_n675), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n682), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n490), .A2(new_n495), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n942), .A2(new_n946), .B1(new_n571), .B2(new_n570), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT111), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n675), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n944), .A2(KEYINPUT42), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n675), .A2(new_n635), .A3(new_n636), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n715), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n624), .A2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n945), .A2(new_n951), .A3(new_n958), .A4(new_n957), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n692), .A2(new_n942), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n699), .B(KEYINPUT41), .Z(new_n967));
  AND3_X1   g0767(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT44), .B1(new_n684), .B2(new_n943), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n682), .A2(new_n683), .A3(new_n942), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT45), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n692), .ZN(new_n974));
  INV_X1    g0774(.A(new_n742), .ZN(new_n975));
  INV_X1    g0775(.A(new_n692), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n685), .B1(new_n529), .B2(new_n675), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n682), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(KEYINPUT112), .B2(new_n691), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n691), .B(KEYINPUT112), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n682), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n967), .B1(new_n985), .B2(new_n975), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n761), .B(KEYINPUT113), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n966), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n229), .A2(new_n755), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n753), .B1(new_n698), .B2(new_n600), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n764), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n826), .A2(new_n472), .B1(new_n798), .B2(new_n447), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G311), .B2(new_n770), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  INV_X1    g0794(.A(G283), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n245), .B1(new_n775), .B2(new_n994), .C1(new_n995), .C2(new_n767), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n786), .B2(G303), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n811), .A2(G116), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n807), .A2(G97), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n993), .A2(new_n997), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n771), .A2(new_n827), .B1(new_n391), .B2(new_n773), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n785), .A2(new_n284), .ZN(new_n1003));
  INV_X1    g0803(.A(G159), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n826), .A2(new_n1004), .B1(new_n798), .B2(new_n214), .ZN(new_n1005));
  INV_X1    g0805(.A(G137), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n254), .B1(new_n775), .B2(new_n1006), .C1(new_n296), .C2(new_n767), .ZN(new_n1007));
  OR4_X1    g0807(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n792), .A2(new_n318), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT47), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n748), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n991), .B1(new_n1012), .B2(new_n1013), .C1(new_n956), .C2(new_n816), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT114), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n983), .A2(new_n742), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n980), .A2(new_n975), .A3(new_n982), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n699), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n773), .A2(new_n318), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1004), .A2(new_n771), .B1(new_n826), .B2(new_n281), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n600), .C2(new_n797), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n254), .B1(new_n775), .B2(new_n284), .C1(new_n214), .C2(new_n767), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n786), .B2(G50), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1000), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(G322), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n826), .A2(new_n804), .B1(new_n771), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT117), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT117), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n786), .A2(G317), .B1(G303), .B2(new_n824), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n798), .A2(new_n995), .B1(new_n773), .B2(new_n472), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n254), .B1(new_n776), .B2(G326), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n514), .C2(new_n792), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT49), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1026), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n748), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n696), .A2(new_n758), .B1(new_n447), .B2(new_n698), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT115), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n696), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n267), .C1(new_n214), .C2(new_n318), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n281), .A2(G50), .ZN(new_n1047));
  XOR2_X1   g0847(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n754), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n233), .A2(new_n267), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n764), .B1(new_n1052), .B2(new_n752), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n685), .B2(new_n751), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n984), .B2(new_n987), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1020), .A2(new_n1056), .ZN(G393));
  INV_X1    g0857(.A(new_n977), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n976), .B1(new_n970), .B2(new_n972), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n987), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n943), .A2(new_n751), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n752), .B1(new_n536), .B2(new_n204), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n241), .A2(new_n755), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n763), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n785), .A2(new_n804), .B1(new_n994), .B2(new_n771), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n245), .B1(new_n767), .B2(new_n472), .C1(new_n798), .C2(new_n514), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1068), .B(new_n793), .C1(G303), .C2(new_n800), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n773), .A2(new_n995), .B1(new_n775), .B2(new_n1027), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT118), .Z(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n785), .A2(new_n1004), .B1(new_n284), .B2(new_n771), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  OAI221_X1 g0874(.A(new_n254), .B1(new_n775), .B2(new_n827), .C1(new_n281), .C2(new_n767), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n798), .A2(new_n318), .B1(new_n773), .B2(new_n214), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G50), .C2(new_n800), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n216), .B2(new_n792), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1065), .B1(new_n1079), .B2(new_n748), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1061), .B1(new_n1062), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1019), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n985), .A3(new_n699), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(G390));
  OAI211_X1 g0884(.A(new_n856), .B(new_n924), .C1(new_n664), .C2(new_n665), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n851), .A2(new_n917), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n885), .A2(new_n887), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n741), .B2(new_n845), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n884), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n843), .A2(new_n372), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n719), .A2(new_n674), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n883), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1087), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1086), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n910), .A2(new_n911), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n889), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n906), .A2(new_n907), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1088), .B1(new_n883), .B2(new_n1093), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n894), .B2(new_n905), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT119), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1094), .A2(new_n888), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n903), .A2(new_n904), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n879), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n912), .B1(new_n1109), .B2(new_n881), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1106), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1102), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT120), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1107), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(KEYINPUT120), .A3(new_n1102), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1087), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1087), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1098), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1117), .A2(KEYINPUT120), .A3(new_n1102), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT120), .B1(new_n1117), .B2(new_n1102), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1121), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1085), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n699), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n764), .B1(new_n838), .B2(new_n281), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT121), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n908), .A2(new_n750), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n826), .A2(new_n447), .B1(new_n771), .B2(new_n995), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n798), .A2(new_n318), .B1(new_n773), .B2(new_n216), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n807), .A2(G68), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n786), .A2(G116), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n245), .B1(new_n775), .B2(new_n472), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G97), .B2(new_n824), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n798), .A2(new_n1004), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n245), .B(new_n1141), .C1(G125), .C2(new_n776), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G128), .A2(new_n770), .B1(new_n800), .B2(G137), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT122), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n824), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n786), .A2(G132), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1142), .A2(new_n1143), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n773), .A2(new_n284), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n296), .B2(new_n792), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1140), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1131), .B(new_n1132), .C1(new_n748), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1121), .B1(new_n1154), .B2(new_n1120), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n987), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1129), .A2(new_n1156), .ZN(G378));
  NAND2_X1  g0957(.A1(new_n301), .A2(new_n673), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n312), .B(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n922), .A2(G330), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n922), .B2(G330), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n914), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n923), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n915), .A3(new_n1163), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n749), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n763), .B1(new_n839), .B2(G50), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n254), .A2(G41), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G50), .B(new_n1173), .C1(new_n251), .C2(new_n266), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1173), .B1(new_n995), .B2(new_n775), .C1(new_n367), .C2(new_n767), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n786), .B2(G107), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n807), .A2(G58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1021), .B1(G68), .B2(new_n797), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G97), .A2(new_n800), .B1(new_n770), .B2(G116), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n786), .A2(G128), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G150), .A2(new_n797), .B1(new_n824), .B2(G137), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G125), .A2(new_n770), .B1(new_n800), .B2(G132), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1145), .A2(new_n811), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1004), .C2(new_n792), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1172), .B1(new_n1192), .B2(new_n748), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1170), .A2(new_n987), .B1(new_n1171), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1085), .B1(new_n1155), .B2(new_n1097), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1164), .A2(new_n1165), .A3(new_n914), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n915), .B1(new_n1168), .B2(new_n1163), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n699), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1128), .A2(new_n1086), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1170), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1199), .B2(new_n1201), .ZN(G375));
  NAND2_X1  g1002(.A1(new_n1088), .A2(new_n749), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n763), .B1(new_n839), .B2(G68), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n771), .A2(new_n472), .B1(new_n798), .B2(new_n367), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n785), .A2(new_n995), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n826), .A2(new_n514), .B1(new_n536), .B2(new_n773), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n254), .B1(new_n776), .B2(G303), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n447), .B2(new_n767), .ZN(new_n1209));
  OR4_X1    g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n767), .A2(new_n284), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n245), .B(new_n1211), .C1(G128), .C2(new_n776), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1145), .A2(new_n800), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n1006), .C2(new_n785), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n770), .A2(G132), .B1(new_n797), .B2(G50), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1177), .B(new_n1215), .C1(new_n1004), .C2(new_n773), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1210), .A2(new_n1009), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1204), .B1(new_n1217), .B2(new_n748), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1203), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1060), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(KEYINPUT123), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1087), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1087), .A2(new_n1089), .B1(new_n883), .B2(new_n848), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n987), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT124), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1224), .A2(new_n1225), .B1(new_n1203), .B2(new_n1218), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT124), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1220), .A2(KEYINPUT123), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n967), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1085), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1098), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G381));
  INV_X1    g1040(.A(G396), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1020), .A2(new_n1056), .A3(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(G390), .A2(G384), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G387), .A2(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(G375), .B(KEYINPUT127), .Z(new_n1246));
  NAND2_X1  g1046(.A1(G378), .A2(KEYINPUT126), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1129), .A2(new_n1248), .A3(new_n1156), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1245), .A2(new_n1246), .A3(new_n1250), .ZN(G407));
  INV_X1    g1051(.A(G343), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G213), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1246), .A2(new_n1250), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  AND2_X1   g1056(.A1(new_n988), .A2(new_n1014), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1242), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1016), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1081), .A2(new_n1083), .B1(new_n1242), .B2(new_n1258), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1257), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1262), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1015), .A3(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1200), .A2(new_n1233), .A3(new_n1170), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1194), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1247), .A2(new_n1249), .A3(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1194), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1253), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(G2897), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1234), .B1(new_n1127), .B2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1085), .A2(new_n1091), .A3(KEYINPUT60), .A4(new_n1096), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n699), .A3(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1221), .A2(new_n1226), .A3(KEYINPUT124), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1229), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G384), .B(new_n1279), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1232), .B2(new_n1279), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n853), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1282), .A3(new_n1274), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1273), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1254), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1267), .A2(new_n1290), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1295), .A2(new_n1298), .A3(new_n1292), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1295), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1295), .B2(new_n1292), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1299), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1297), .B1(new_n1304), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1105(.A1(new_n1250), .A2(G375), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1293), .A3(new_n1271), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1293), .B1(new_n1306), .B2(new_n1271), .ZN(new_n1310));
  OR3_X1    g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


