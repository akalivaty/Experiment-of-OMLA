

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783;

  AND2_X1 U376 ( .A1(n427), .A2(n426), .ZN(n430) );
  NAND2_X1 U377 ( .A1(n451), .A2(n456), .ZN(n601) );
  INV_X1 U378 ( .A(n706), .ZN(n456) );
  NOR2_X1 U379 ( .A1(n707), .A2(n706), .ZN(n649) );
  XNOR2_X1 U380 ( .A(n391), .B(n522), .ZN(n574) );
  INV_X1 U381 ( .A(G953), .ZN(n769) );
  AND2_X4 U382 ( .A1(n389), .A2(n699), .ZN(n744) );
  OR2_X2 U383 ( .A1(n746), .A2(G902), .ZN(n531) );
  XNOR2_X2 U384 ( .A(n629), .B(KEYINPUT22), .ZN(n635) );
  XNOR2_X2 U385 ( .A(n575), .B(n753), .ZN(n742) );
  XNOR2_X1 U386 ( .A(n649), .B(KEYINPUT105), .ZN(n431) );
  INV_X4 U387 ( .A(G143), .ZN(n483) );
  NAND2_X1 U388 ( .A1(n387), .A2(n386), .ZN(n389) );
  XNOR2_X1 U389 ( .A(n662), .B(KEYINPUT103), .ZN(n663) );
  XNOR2_X1 U390 ( .A(n493), .B(n492), .ZN(n781) );
  NAND2_X1 U391 ( .A1(n371), .A2(n384), .ZN(n379) );
  XNOR2_X1 U392 ( .A(n590), .B(KEYINPUT1), .ZN(n707) );
  OR2_X2 U393 ( .A1(n517), .A2(n604), .ZN(n689) );
  XNOR2_X1 U394 ( .A(n418), .B(n504), .ZN(n669) );
  XNOR2_X1 U395 ( .A(n458), .B(n457), .ZN(n523) );
  NOR2_X1 U396 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n639) );
  BUF_X1 U397 ( .A(n624), .Z(n357) );
  XNOR2_X1 U398 ( .A(n428), .B(KEYINPUT104), .ZN(n358) );
  XNOR2_X1 U399 ( .A(n370), .B(KEYINPUT19), .ZN(n624) );
  XNOR2_X1 U400 ( .A(n428), .B(KEYINPUT104), .ZN(n779) );
  XNOR2_X1 U401 ( .A(n468), .B(n467), .ZN(n370) );
  XNOR2_X2 U402 ( .A(n645), .B(n644), .ZN(n777) );
  XNOR2_X1 U403 ( .A(n570), .B(n482), .ZN(n524) );
  XNOR2_X2 U404 ( .A(n573), .B(n412), .ZN(n440) );
  NOR2_X2 U405 ( .A1(n614), .A2(n579), .ZN(n468) );
  NOR2_X1 U406 ( .A1(n588), .A2(n780), .ZN(n589) );
  XNOR2_X1 U407 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n509) );
  XNOR2_X1 U408 ( .A(n525), .B(n523), .ZN(n538) );
  XNOR2_X1 U409 ( .A(n524), .B(KEYINPUT69), .ZN(n525) );
  AND2_X1 U410 ( .A1(n592), .A2(n489), .ZN(n486) );
  XNOR2_X1 U411 ( .A(n576), .B(KEYINPUT89), .ZN(n577) );
  NAND2_X1 U412 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U413 ( .A(n379), .ZN(n383) );
  XOR2_X1 U414 ( .A(KEYINPUT87), .B(G110), .Z(n522) );
  XNOR2_X1 U415 ( .A(n521), .B(n439), .ZN(n391) );
  INV_X1 U416 ( .A(G107), .ZN(n439) );
  XNOR2_X1 U417 ( .A(n538), .B(n495), .ZN(n765) );
  INV_X1 U418 ( .A(n547), .ZN(n495) );
  XNOR2_X1 U419 ( .A(n400), .B(G101), .ZN(n565) );
  INV_X1 U420 ( .A(KEYINPUT4), .ZN(n400) );
  INV_X1 U421 ( .A(KEYINPUT108), .ZN(n441) );
  NAND2_X1 U422 ( .A1(n603), .A2(n491), .ZN(n489) );
  XNOR2_X1 U423 ( .A(n515), .B(G478), .ZN(n604) );
  INV_X1 U424 ( .A(KEYINPUT66), .ZN(n457) );
  XNOR2_X1 U425 ( .A(G131), .B(KEYINPUT67), .ZN(n458) );
  XNOR2_X1 U426 ( .A(n477), .B(n476), .ZN(n459) );
  OR2_X1 U427 ( .A1(G902), .A2(G237), .ZN(n578) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n532) );
  XNOR2_X1 U429 ( .A(G137), .B(KEYINPUT68), .ZN(n547) );
  XNOR2_X1 U430 ( .A(n506), .B(G475), .ZN(n465) );
  OR2_X1 U431 ( .A1(n669), .A2(G902), .ZN(n466) );
  XNOR2_X1 U432 ( .A(n704), .B(KEYINPUT6), .ZN(n641) );
  XNOR2_X1 U433 ( .A(n569), .B(n442), .ZN(n764) );
  XNOR2_X1 U434 ( .A(n526), .B(KEYINPUT10), .ZN(n442) );
  XNOR2_X1 U435 ( .A(G128), .B(G110), .ZN(n543) );
  XNOR2_X1 U436 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n496) );
  XNOR2_X1 U437 ( .A(n566), .B(n473), .ZN(n472) );
  INV_X1 U438 ( .A(KEYINPUT18), .ZN(n473) );
  XNOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT88), .ZN(n566) );
  OR2_X1 U440 ( .A1(n432), .A2(n364), .ZN(n394) );
  AND2_X1 U441 ( .A1(n432), .A2(n364), .ZN(n396) );
  XNOR2_X1 U442 ( .A(n689), .B(n516), .ZN(n616) );
  INV_X1 U443 ( .A(KEYINPUT99), .ZN(n516) );
  AND2_X1 U444 ( .A1(n486), .A2(n456), .ZN(n409) );
  NAND2_X1 U445 ( .A1(n484), .A2(n362), .ZN(n487) );
  AND2_X1 U446 ( .A1(n378), .A2(n376), .ZN(n375) );
  NAND2_X1 U447 ( .A1(n379), .A2(n385), .ZN(n378) );
  NAND2_X1 U448 ( .A1(n377), .A2(n385), .ZN(n376) );
  NAND2_X1 U449 ( .A1(n380), .A2(KEYINPUT34), .ZN(n374) );
  BUF_X1 U450 ( .A(n707), .Z(n432) );
  AND2_X1 U451 ( .A1(n452), .A2(n453), .ZN(n451) );
  AND2_X1 U452 ( .A1(n455), .A2(n584), .ZN(n452) );
  XNOR2_X1 U453 ( .A(n583), .B(n454), .ZN(n453) );
  INV_X1 U454 ( .A(KEYINPUT30), .ZN(n454) );
  AND2_X1 U455 ( .A1(n456), .A2(n449), .ZN(n450) );
  OR2_X1 U456 ( .A1(n749), .A2(G902), .ZN(n448) );
  XOR2_X1 U457 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n555) );
  XNOR2_X1 U458 ( .A(n671), .B(n368), .ZN(n672) );
  XNOR2_X1 U459 ( .A(n413), .B(G122), .ZN(n412) );
  XNOR2_X1 U460 ( .A(KEYINPUT16), .B(KEYINPUT70), .ZN(n413) );
  NAND2_X1 U461 ( .A1(n666), .A2(KEYINPUT2), .ZN(n386) );
  NAND2_X1 U462 ( .A1(n417), .A2(n359), .ZN(n387) );
  XNOR2_X1 U463 ( .A(n513), .B(n437), .ZN(n747) );
  XNOR2_X1 U464 ( .A(n670), .B(n471), .ZN(n470) );
  INV_X1 U465 ( .A(KEYINPUT59), .ZN(n471) );
  XNOR2_X1 U466 ( .A(n529), .B(n528), .ZN(n494) );
  XNOR2_X1 U467 ( .A(n527), .B(n526), .ZN(n528) );
  NOR2_X1 U468 ( .A1(n402), .A2(n401), .ZN(n478) );
  INV_X1 U469 ( .A(KEYINPUT72), .ZN(n535) );
  XNOR2_X1 U470 ( .A(G137), .B(KEYINPUT5), .ZN(n536) );
  XNOR2_X1 U471 ( .A(n408), .B(KEYINPUT81), .ZN(n416) );
  XNOR2_X1 U472 ( .A(G902), .B(KEYINPUT15), .ZN(n540) );
  XNOR2_X1 U473 ( .A(G104), .B(KEYINPUT73), .ZN(n521) );
  XNOR2_X1 U474 ( .A(KEYINPUT65), .B(n582), .ZN(n706) );
  INV_X1 U475 ( .A(n416), .ZN(n767) );
  XOR2_X1 U476 ( .A(KEYINPUT98), .B(G122), .Z(n508) );
  XNOR2_X1 U477 ( .A(G107), .B(G116), .ZN(n507) );
  XOR2_X1 U478 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n512) );
  INV_X1 U479 ( .A(G134), .ZN(n482) );
  XNOR2_X1 U480 ( .A(n505), .B(n764), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n565), .B(n399), .ZN(n534) );
  INV_X1 U482 ( .A(G146), .ZN(n399) );
  NOR2_X1 U483 ( .A1(n593), .A2(n641), .ZN(n594) );
  INV_X1 U484 ( .A(KEYINPUT84), .ZN(n467) );
  XNOR2_X1 U485 ( .A(n605), .B(KEYINPUT97), .ZN(n517) );
  OR2_X1 U486 ( .A1(n671), .A2(G902), .ZN(n398) );
  INV_X1 U487 ( .A(n590), .ZN(n455) );
  INV_X1 U488 ( .A(n641), .ZN(n657) );
  XNOR2_X1 U489 ( .A(n551), .B(n552), .ZN(n749) );
  XNOR2_X1 U490 ( .A(n764), .B(n546), .ZN(n552) );
  XNOR2_X1 U491 ( .A(n545), .B(n496), .ZN(n546) );
  XNOR2_X1 U492 ( .A(n429), .B(n568), .ZN(n575) );
  XNOR2_X1 U493 ( .A(n472), .B(n565), .ZN(n568) );
  XNOR2_X1 U494 ( .A(n572), .B(n567), .ZN(n429) );
  NAND2_X1 U495 ( .A1(n393), .A2(n392), .ZN(n694) );
  AND2_X1 U496 ( .A1(n395), .A2(n363), .ZN(n393) );
  NAND2_X1 U497 ( .A1(n488), .A2(n487), .ZN(n615) );
  INV_X1 U498 ( .A(KEYINPUT40), .ZN(n492) );
  NAND2_X1 U499 ( .A1(n411), .A2(n410), .ZN(n485) );
  NAND2_X1 U500 ( .A1(n375), .A2(n372), .ZN(n643) );
  NAND2_X1 U501 ( .A1(n450), .A2(n451), .ZN(n586) );
  INV_X1 U502 ( .A(KEYINPUT63), .ZN(n433) );
  XNOR2_X1 U503 ( .A(n481), .B(n480), .ZN(n479) );
  INV_X1 U504 ( .A(n747), .ZN(n480) );
  XNOR2_X1 U505 ( .A(n668), .B(n470), .ZN(n469) );
  NAND2_X1 U506 ( .A1(n463), .A2(n426), .ZN(n462) );
  XNOR2_X1 U507 ( .A(n464), .B(n366), .ZN(n463) );
  XNOR2_X1 U508 ( .A(n740), .B(n422), .ZN(G75) );
  XNOR2_X1 U509 ( .A(n423), .B(KEYINPUT53), .ZN(n422) );
  INV_X1 U510 ( .A(KEYINPUT120), .ZN(n423) );
  AND2_X1 U511 ( .A1(n416), .A2(n666), .ZN(n359) );
  AND2_X1 U512 ( .A1(n456), .A2(n455), .ZN(n360) );
  OR2_X1 U513 ( .A1(n683), .A2(n599), .ZN(n361) );
  BUF_X1 U514 ( .A(n614), .Z(n438) );
  INV_X1 U515 ( .A(n438), .ZN(n449) );
  NOR2_X1 U516 ( .A1(n603), .A2(n491), .ZN(n362) );
  INV_X1 U517 ( .A(G140), .ZN(n526) );
  AND2_X1 U518 ( .A1(n394), .A2(n438), .ZN(n363) );
  XOR2_X1 U519 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n364) );
  XOR2_X1 U520 ( .A(KEYINPUT33), .B(KEYINPUT106), .Z(n365) );
  INV_X1 U521 ( .A(KEYINPUT39), .ZN(n491) );
  XOR2_X1 U522 ( .A(n746), .B(n745), .Z(n366) );
  XOR2_X1 U523 ( .A(n742), .B(n741), .Z(n367) );
  INV_X1 U524 ( .A(KEYINPUT34), .ZN(n385) );
  NOR2_X1 U525 ( .A1(G952), .A2(n769), .ZN(n750) );
  INV_X1 U526 ( .A(n750), .ZN(n426) );
  XNOR2_X1 U527 ( .A(KEYINPUT62), .B(KEYINPUT86), .ZN(n368) );
  XOR2_X1 U528 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n369) );
  NOR2_X1 U529 ( .A1(n611), .A2(n370), .ZN(n595) );
  NAND2_X1 U530 ( .A1(n431), .A2(n365), .ZN(n371) );
  NAND2_X1 U531 ( .A1(n383), .A2(n380), .ZN(n734) );
  NAND2_X1 U532 ( .A1(n373), .A2(n383), .ZN(n372) );
  NOR2_X1 U533 ( .A1(n374), .A2(n650), .ZN(n373) );
  NAND2_X1 U534 ( .A1(n652), .A2(n380), .ZN(n377) );
  NOR2_X1 U535 ( .A1(n641), .A2(n365), .ZN(n381) );
  INV_X1 U536 ( .A(n431), .ZN(n382) );
  NAND2_X1 U537 ( .A1(n641), .A2(n365), .ZN(n384) );
  XNOR2_X2 U538 ( .A(n388), .B(KEYINPUT74), .ZN(n699) );
  NAND2_X1 U539 ( .A1(n667), .A2(n474), .ZN(n388) );
  XNOR2_X2 U540 ( .A(n665), .B(KEYINPUT45), .ZN(n667) );
  INV_X2 U541 ( .A(G125), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n390), .B(n523), .ZN(n505) );
  XNOR2_X1 U543 ( .A(n499), .B(n498), .ZN(n390) );
  NAND2_X1 U544 ( .A1(n459), .A2(n618), .ZN(n408) );
  OR2_X1 U545 ( .A1(n397), .A2(n364), .ZN(n392) );
  NAND2_X1 U546 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U547 ( .A(n613), .B(n441), .ZN(n397) );
  XNOR2_X2 U548 ( .A(n398), .B(G472), .ZN(n704) );
  NAND2_X1 U549 ( .A1(n361), .A2(n403), .ZN(n401) );
  NAND2_X1 U550 ( .A1(n405), .A2(n404), .ZN(n402) );
  NAND2_X1 U551 ( .A1(n782), .A2(KEYINPUT46), .ZN(n403) );
  NAND2_X1 U552 ( .A1(n781), .A2(KEYINPUT46), .ZN(n404) );
  NAND2_X1 U553 ( .A1(n407), .A2(n406), .ZN(n405) );
  NOR2_X1 U554 ( .A1(n782), .A2(KEYINPUT46), .ZN(n406) );
  INV_X1 U555 ( .A(n781), .ZN(n407) );
  NAND2_X1 U556 ( .A1(n409), .A2(n451), .ZN(n411) );
  NAND2_X1 U557 ( .A1(n601), .A2(n491), .ZN(n490) );
  NAND2_X1 U558 ( .A1(n486), .A2(KEYINPUT39), .ZN(n410) );
  XNOR2_X2 U559 ( .A(n415), .B(n414), .ZN(n573) );
  XNOR2_X2 U560 ( .A(G119), .B(G116), .ZN(n414) );
  XNOR2_X2 U561 ( .A(n435), .B(G113), .ZN(n415) );
  INV_X1 U562 ( .A(n759), .ZN(n417) );
  INV_X1 U563 ( .A(KEYINPUT44), .ZN(n419) );
  XNOR2_X1 U564 ( .A(n765), .B(n494), .ZN(n746) );
  NAND2_X1 U565 ( .A1(n659), .A2(n632), .ZN(n428) );
  NAND2_X1 U566 ( .A1(n744), .A2(G217), .ZN(n748) );
  INV_X2 U567 ( .A(KEYINPUT3), .ZN(n435) );
  NAND2_X1 U568 ( .A1(n420), .A2(n419), .ZN(n647) );
  INV_X1 U569 ( .A(n777), .ZN(n420) );
  NOR2_X2 U570 ( .A1(n742), .A2(n666), .ZN(n421) );
  XNOR2_X2 U571 ( .A(n421), .B(n577), .ZN(n614) );
  XNOR2_X1 U572 ( .A(n461), .B(n475), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n424), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U574 ( .A1(n479), .A2(n426), .ZN(n424) );
  XNOR2_X1 U575 ( .A(n425), .B(n369), .ZN(G60) );
  NAND2_X1 U576 ( .A1(n469), .A2(n426), .ZN(n425) );
  XNOR2_X1 U577 ( .A(n743), .B(n367), .ZN(n427) );
  NAND2_X1 U578 ( .A1(n485), .A2(n487), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n430), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U580 ( .A(n434), .B(n433), .ZN(G57) );
  NOR2_X2 U581 ( .A1(n674), .A2(n750), .ZN(n434) );
  XNOR2_X1 U582 ( .A(n436), .B(n533), .ZN(n539) );
  XNOR2_X1 U583 ( .A(n534), .B(n537), .ZN(n436) );
  XNOR2_X1 U584 ( .A(n524), .B(n514), .ZN(n437) );
  NAND2_X1 U585 ( .A1(n779), .A2(n778), .ZN(n640) );
  XNOR2_X2 U586 ( .A(n638), .B(KEYINPUT32), .ZN(n778) );
  XNOR2_X2 U587 ( .A(n440), .B(n574), .ZN(n753) );
  XNOR2_X1 U588 ( .A(n594), .B(KEYINPUT107), .ZN(n611) );
  XNOR2_X2 U589 ( .A(n443), .B(G146), .ZN(n569) );
  NAND2_X1 U590 ( .A1(n444), .A2(n739), .ZN(n740) );
  NAND2_X1 U591 ( .A1(n445), .A2(n699), .ZN(n444) );
  XNOR2_X1 U592 ( .A(n447), .B(n446), .ZN(n445) );
  INV_X1 U593 ( .A(KEYINPUT76), .ZN(n446) );
  NAND2_X1 U594 ( .A1(n698), .A2(n697), .ZN(n447) );
  NOR2_X1 U595 ( .A1(n633), .A2(n701), .ZN(n582) );
  XNOR2_X2 U596 ( .A(n448), .B(n556), .ZN(n633) );
  NAND2_X1 U597 ( .A1(n767), .A2(n696), .ZN(n695) );
  NAND2_X1 U598 ( .A1(n460), .A2(n459), .ZN(n461) );
  AND2_X1 U599 ( .A1(n618), .A2(KEYINPUT2), .ZN(n460) );
  XNOR2_X1 U600 ( .A(n462), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U601 ( .A1(n744), .A2(G469), .ZN(n464) );
  XNOR2_X2 U602 ( .A(n466), .B(n465), .ZN(n605) );
  NAND2_X1 U603 ( .A1(n624), .A2(n623), .ZN(n627) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U605 ( .A(n611), .ZN(n612) );
  INV_X1 U606 ( .A(KEYINPUT82), .ZN(n475) );
  INV_X1 U607 ( .A(KEYINPUT48), .ZN(n476) );
  NAND2_X1 U608 ( .A1(n610), .A2(n478), .ZN(n477) );
  NAND2_X1 U609 ( .A1(n744), .A2(G478), .ZN(n481) );
  XNOR2_X2 U610 ( .A(n483), .B(G128), .ZN(n570) );
  INV_X1 U611 ( .A(n601), .ZN(n484) );
  AND2_X1 U612 ( .A1(n490), .A2(n489), .ZN(n488) );
  NOR2_X2 U613 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U614 ( .A1(G210), .A2(n532), .ZN(n497) );
  INV_X1 U615 ( .A(KEYINPUT100), .ZN(n518) );
  XNOR2_X1 U616 ( .A(n536), .B(n535), .ZN(n537) );
  INV_X1 U617 ( .A(n571), .ZN(n572) );
  INV_X1 U618 ( .A(G469), .ZN(n530) );
  INV_X1 U619 ( .A(n669), .ZN(n670) );
  XNOR2_X1 U620 ( .A(n673), .B(n672), .ZN(n674) );
  INV_X1 U621 ( .A(n540), .ZN(n666) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n499) );
  XNOR2_X1 U623 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n498) );
  XOR2_X1 U624 ( .A(G113), .B(G104), .Z(n501) );
  XNOR2_X1 U625 ( .A(G143), .B(G122), .ZN(n500) );
  XNOR2_X1 U626 ( .A(n500), .B(n501), .ZN(n503) );
  NAND2_X1 U627 ( .A1(n532), .A2(G214), .ZN(n502) );
  XNOR2_X1 U628 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n506) );
  XNOR2_X1 U629 ( .A(n508), .B(n507), .ZN(n514) );
  NAND2_X1 U630 ( .A1(n769), .A2(G234), .ZN(n510) );
  XNOR2_X1 U631 ( .A(n510), .B(n509), .ZN(n548) );
  NAND2_X1 U632 ( .A1(G217), .A2(n548), .ZN(n511) );
  XNOR2_X1 U633 ( .A(n512), .B(n511), .ZN(n513) );
  NOR2_X1 U634 ( .A1(G902), .A2(n747), .ZN(n515) );
  NAND2_X1 U635 ( .A1(n604), .A2(n517), .ZN(n685) );
  NAND2_X1 U636 ( .A1(n616), .A2(n685), .ZN(n519) );
  XNOR2_X2 U637 ( .A(n519), .B(n518), .ZN(n723) );
  NAND2_X1 U638 ( .A1(n723), .A2(KEYINPUT47), .ZN(n520) );
  XNOR2_X1 U639 ( .A(n520), .B(KEYINPUT78), .ZN(n581) );
  XNOR2_X1 U640 ( .A(n574), .B(n534), .ZN(n529) );
  NAND2_X1 U641 ( .A1(G227), .A2(n769), .ZN(n527) );
  XNOR2_X2 U642 ( .A(n531), .B(n530), .ZN(n590) );
  XNOR2_X1 U643 ( .A(n573), .B(n497), .ZN(n533) );
  XNOR2_X1 U644 ( .A(n538), .B(n539), .ZN(n671) );
  NAND2_X1 U645 ( .A1(G234), .A2(n540), .ZN(n541) );
  XNOR2_X1 U646 ( .A(KEYINPUT20), .B(n541), .ZN(n553) );
  NAND2_X1 U647 ( .A1(G221), .A2(n553), .ZN(n542) );
  XNOR2_X1 U648 ( .A(n542), .B(KEYINPUT21), .ZN(n701) );
  XOR2_X1 U649 ( .A(KEYINPUT23), .B(G119), .Z(n544) );
  XNOR2_X1 U650 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U651 ( .A(n547), .B(KEYINPUT24), .ZN(n550) );
  NAND2_X1 U652 ( .A1(G221), .A2(n548), .ZN(n549) );
  XNOR2_X1 U653 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U654 ( .A1(n553), .A2(G217), .ZN(n554) );
  XNOR2_X1 U655 ( .A(n555), .B(n554), .ZN(n556) );
  NAND2_X1 U656 ( .A1(G237), .A2(G234), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n557), .B(KEYINPUT14), .ZN(n559) );
  NAND2_X1 U658 ( .A1(G952), .A2(n559), .ZN(n732) );
  NOR2_X1 U659 ( .A1(G953), .A2(n732), .ZN(n558) );
  XOR2_X1 U660 ( .A(KEYINPUT90), .B(n558), .Z(n621) );
  NAND2_X1 U661 ( .A1(G902), .A2(n559), .ZN(n619) );
  NOR2_X1 U662 ( .A1(G900), .A2(n619), .ZN(n560) );
  NAND2_X1 U663 ( .A1(G953), .A2(n560), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n621), .A2(n561), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n633), .A2(n584), .ZN(n562) );
  NOR2_X1 U666 ( .A1(n701), .A2(n562), .ZN(n591) );
  AND2_X1 U667 ( .A1(n704), .A2(n591), .ZN(n563) );
  XOR2_X1 U668 ( .A(KEYINPUT28), .B(n563), .Z(n564) );
  NOR2_X1 U669 ( .A1(n590), .A2(n564), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G224), .A2(n769), .ZN(n567) );
  XNOR2_X1 U671 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U672 ( .A1(G210), .A2(n578), .ZN(n576) );
  NAND2_X1 U673 ( .A1(G214), .A2(n578), .ZN(n718) );
  INV_X1 U674 ( .A(n718), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n602), .A2(n357), .ZN(n683) );
  NAND2_X1 U676 ( .A1(n683), .A2(KEYINPUT47), .ZN(n580) );
  NAND2_X1 U677 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n704), .A2(n718), .ZN(n583) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n642) );
  INV_X1 U680 ( .A(n642), .ZN(n585) );
  NOR2_X1 U681 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U682 ( .A(n587), .B(KEYINPUT110), .ZN(n780) );
  XNOR2_X1 U683 ( .A(KEYINPUT77), .B(n589), .ZN(n597) );
  INV_X1 U684 ( .A(n685), .ZN(n592) );
  NAND2_X1 U685 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U686 ( .A(KEYINPUT36), .B(n595), .Z(n596) );
  NOR2_X1 U687 ( .A1(n432), .A2(n596), .ZN(n691) );
  NOR2_X1 U688 ( .A1(n597), .A2(n691), .ZN(n610) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n723), .ZN(n598) );
  XNOR2_X1 U690 ( .A(n598), .B(KEYINPUT71), .ZN(n599) );
  INV_X1 U691 ( .A(KEYINPUT38), .ZN(n600) );
  XNOR2_X1 U692 ( .A(n614), .B(n600), .ZN(n603) );
  INV_X1 U693 ( .A(n602), .ZN(n607) );
  INV_X1 U694 ( .A(n603), .ZN(n719) );
  NAND2_X1 U695 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U696 ( .A1(n605), .A2(n604), .ZN(n722) );
  NOR2_X1 U697 ( .A1(n724), .A2(n722), .ZN(n606) );
  XNOR2_X1 U698 ( .A(n606), .B(KEYINPUT41), .ZN(n733) );
  NOR2_X1 U699 ( .A1(n607), .A2(n733), .ZN(n609) );
  XOR2_X1 U700 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n608) );
  XNOR2_X1 U701 ( .A(n609), .B(n608), .ZN(n782) );
  NAND2_X1 U702 ( .A1(n612), .A2(n718), .ZN(n613) );
  NOR2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n693) );
  INV_X1 U704 ( .A(n693), .ZN(n617) );
  AND2_X1 U705 ( .A1(n694), .A2(n617), .ZN(n618) );
  NOR2_X1 U706 ( .A1(G898), .A2(n769), .ZN(n755) );
  INV_X1 U707 ( .A(n619), .ZN(n620) );
  NAND2_X1 U708 ( .A1(n755), .A2(n620), .ZN(n622) );
  NAND2_X1 U709 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U710 ( .A(KEYINPUT0), .B(KEYINPUT64), .ZN(n625) );
  XNOR2_X1 U711 ( .A(n625), .B(KEYINPUT85), .ZN(n626) );
  XNOR2_X2 U712 ( .A(n627), .B(n626), .ZN(n652) );
  NOR2_X1 U713 ( .A1(n701), .A2(n722), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n652), .A2(n628), .ZN(n629) );
  INV_X1 U715 ( .A(n432), .ZN(n630) );
  NOR2_X2 U716 ( .A1(n635), .A2(n630), .ZN(n659) );
  INV_X1 U717 ( .A(n633), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n631), .A2(n704), .ZN(n632) );
  XOR2_X1 U719 ( .A(KEYINPUT101), .B(n633), .Z(n700) );
  INV_X1 U720 ( .A(n700), .ZN(n634) );
  NOR2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n657), .A2(n432), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U724 ( .A(n640), .B(n639), .ZN(n646) );
  INV_X1 U725 ( .A(n652), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  INV_X1 U727 ( .A(KEYINPUT35), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n646), .A2(n777), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n704), .A2(n649), .ZN(n713) );
  NOR2_X1 U731 ( .A1(n713), .A2(n650), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n651), .B(KEYINPUT31), .ZN(n688) );
  NAND2_X1 U733 ( .A1(n652), .A2(n360), .ZN(n653) );
  NOR2_X1 U734 ( .A1(n704), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n654), .B(KEYINPUT93), .ZN(n678) );
  NAND2_X1 U736 ( .A1(n688), .A2(n678), .ZN(n656) );
  INV_X1 U737 ( .A(n723), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n661) );
  NOR2_X1 U739 ( .A1(n657), .A2(n700), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U741 ( .A(KEYINPUT102), .B(n660), .ZN(n783) );
  NAND2_X1 U742 ( .A1(n661), .A2(n783), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(n665) );
  INV_X1 U744 ( .A(n667), .ZN(n759) );
  NAND2_X1 U745 ( .A1(n744), .A2(G475), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n744), .A2(G472), .ZN(n673) );
  NOR2_X1 U747 ( .A1(n685), .A2(n678), .ZN(n675) );
  XOR2_X1 U748 ( .A(G104), .B(n675), .Z(G6) );
  XOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n677) );
  XNOR2_X1 U750 ( .A(G107), .B(KEYINPUT112), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n689), .A2(n678), .ZN(n679) );
  XOR2_X1 U753 ( .A(n680), .B(n679), .Z(G9) );
  NOR2_X1 U754 ( .A1(n689), .A2(n683), .ZN(n682) );
  XNOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .ZN(n681) );
  XNOR2_X1 U756 ( .A(n682), .B(n681), .ZN(G30) );
  NOR2_X1 U757 ( .A1(n685), .A2(n683), .ZN(n684) );
  XOR2_X1 U758 ( .A(G146), .B(n684), .Z(G48) );
  NOR2_X1 U759 ( .A1(n685), .A2(n688), .ZN(n687) );
  XNOR2_X1 U760 ( .A(G113), .B(KEYINPUT113), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(G15) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U763 ( .A(G116), .B(n690), .Z(G18) );
  XNOR2_X1 U764 ( .A(G125), .B(n691), .ZN(n692) );
  XNOR2_X1 U765 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U766 ( .A(G134), .B(n693), .Z(G36) );
  XNOR2_X1 U767 ( .A(n694), .B(G140), .ZN(G42) );
  INV_X1 U768 ( .A(KEYINPUT2), .ZN(n696) );
  XNOR2_X1 U769 ( .A(n695), .B(KEYINPUT80), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n759), .A2(n696), .ZN(n697) );
  NAND2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n702), .ZN(n703) );
  NOR2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U774 ( .A(KEYINPUT114), .B(n705), .ZN(n711) );
  XOR2_X1 U775 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n709) );
  NAND2_X1 U776 ( .A1(n432), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n712), .B(KEYINPUT116), .ZN(n714) );
  NAND2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U781 ( .A(KEYINPUT51), .B(n715), .ZN(n716) );
  NOR2_X1 U782 ( .A1(n733), .A2(n716), .ZN(n717) );
  XOR2_X1 U783 ( .A(KEYINPUT117), .B(n717), .Z(n729) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(n720), .B(KEYINPUT118), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U789 ( .A1(n734), .A2(n727), .ZN(n728) );
  NOR2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U791 ( .A(n730), .B(KEYINPUT52), .ZN(n731) );
  NOR2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n738) );
  NOR2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U794 ( .A(n735), .B(KEYINPUT119), .ZN(n736) );
  NAND2_X1 U795 ( .A1(n769), .A2(n736), .ZN(n737) );
  NOR2_X1 U796 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U797 ( .A1(n744), .A2(G210), .ZN(n743) );
  XOR2_X1 U798 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n741) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  XNOR2_X1 U800 ( .A(n748), .B(n749), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(KEYINPUT124), .ZN(G66) );
  XOR2_X1 U802 ( .A(n753), .B(G101), .Z(n754) );
  NOR2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n763) );
  XOR2_X1 U804 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n757) );
  NAND2_X1 U805 ( .A1(G224), .A2(G953), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G898), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n417), .A2(n769), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U810 ( .A(n763), .B(n762), .ZN(G69) );
  XOR2_X1 U811 ( .A(n764), .B(KEYINPUT4), .Z(n766) );
  XNOR2_X1 U812 ( .A(n766), .B(n765), .ZN(n771) );
  XNOR2_X1 U813 ( .A(KEYINPUT126), .B(n767), .ZN(n768) );
  XNOR2_X1 U814 ( .A(n771), .B(n768), .ZN(n770) );
  NAND2_X1 U815 ( .A1(n770), .A2(n769), .ZN(n776) );
  XNOR2_X1 U816 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U817 ( .A1(n772), .A2(G900), .ZN(n773) );
  XOR2_X1 U818 ( .A(KEYINPUT127), .B(n773), .Z(n774) );
  NAND2_X1 U819 ( .A1(G953), .A2(n774), .ZN(n775) );
  NAND2_X1 U820 ( .A1(n776), .A2(n775), .ZN(G72) );
  XNOR2_X1 U821 ( .A(n777), .B(G122), .ZN(G24) );
  XNOR2_X1 U822 ( .A(n778), .B(G119), .ZN(G21) );
  XNOR2_X1 U823 ( .A(n358), .B(G110), .ZN(G12) );
  XOR2_X1 U824 ( .A(G143), .B(n780), .Z(G45) );
  XOR2_X1 U825 ( .A(n781), .B(G131), .Z(G33) );
  XOR2_X1 U826 ( .A(G137), .B(n782), .Z(G39) );
  XNOR2_X1 U827 ( .A(G101), .B(n783), .ZN(G3) );
endmodule

