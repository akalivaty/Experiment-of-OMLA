//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI22_X1  g001(.A1(new_n187), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(G104), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G104), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n190), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n191), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n202), .B(G146), .C1(new_n203), .C2(KEYINPUT1), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT67), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n211), .A4(G128), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n201), .A2(KEYINPUT10), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n201), .A2(KEYINPUT81), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT81), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n197), .A2(new_n221), .A3(new_n200), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n225), .A3(new_n206), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n220), .A2(new_n222), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n219), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n190), .A2(new_n194), .A3(G101), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n195), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT79), .B1(new_n190), .B2(new_n194), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n233), .A2(new_n234), .A3(G101), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n231), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n235), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(new_n196), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n234), .A3(KEYINPUT4), .A4(new_n233), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n214), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n210), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n230), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n227), .A2(new_n223), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n197), .A2(new_n221), .A3(new_n200), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n221), .B1(new_n197), .B2(new_n200), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n218), .B1(new_n256), .B2(KEYINPUT10), .ZN(new_n257));
  INV_X1    g071(.A(new_n248), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n210), .A2(new_n243), .A3(new_n247), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n238), .B2(new_n241), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT83), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT65), .B(G131), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(new_n265), .A3(new_n267), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n252), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n275), .B(new_n277), .Z(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n257), .A2(new_n261), .ZN(new_n280));
  INV_X1    g094(.A(new_n273), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n230), .A2(new_n250), .A3(new_n281), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n201), .A2(new_n223), .A3(new_n227), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n201), .B2(new_n217), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n286), .A2(KEYINPUT82), .A3(new_n287), .A4(new_n273), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(KEYINPUT82), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n287), .A2(KEYINPUT82), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n284), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT84), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n282), .A2(new_n274), .B1(new_n293), .B2(new_n279), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n298), .B(G469), .C1(new_n299), .C2(G902), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n288), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT85), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n304), .A3(new_n288), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n303), .A2(new_n282), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n278), .B1(new_n274), .B2(new_n284), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n296), .B(new_n301), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n297), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G221), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT9), .B(G234), .Z(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n301), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G116), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n238), .B2(new_n241), .ZN(new_n324));
  XOR2_X1   g138(.A(G110), .B(G122), .Z(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n327));
  INV_X1    g141(.A(G113), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n321), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(new_n322), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n220), .B2(new_n222), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n324), .A2(new_n325), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n325), .B1(new_n324), .B2(new_n333), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n260), .A2(G125), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n253), .B2(G125), .ZN(new_n338));
  INV_X1    g152(.A(G224), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G953), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT86), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(new_n325), .C1(new_n324), .C2(new_n333), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT7), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n338), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n338), .A2(new_n340), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n329), .B1(new_n326), .B2(KEYINPUT87), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(KEYINPUT87), .B2(new_n326), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n331), .A2(new_n322), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n351), .A2(new_n201), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n353), .A2(new_n354), .B1(new_n201), .B2(new_n332), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n201), .A2(new_n352), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT88), .B1(new_n356), .B2(new_n351), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n325), .B(KEYINPUT8), .Z(new_n359));
  AOI21_X1  g173(.A(new_n349), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n360), .B2(new_n334), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n345), .A2(new_n361), .A3(new_n363), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n316), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n276), .A2(G952), .ZN(new_n368));
  NAND2_X1  g182(.A1(G234), .A2(G237), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT21), .B(G898), .Z(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(G902), .A3(G953), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n203), .A2(G143), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n203), .A2(G143), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n264), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT96), .B(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n319), .A2(G122), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n189), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n319), .A3(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT98), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n379), .B(new_n383), .C1(new_n388), .C2(new_n189), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(new_n382), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n383), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT97), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n377), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n393), .A2(KEYINPUT97), .ZN(new_n397));
  OAI21_X1  g211(.A(G134), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n378), .A2(new_n264), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n392), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n311), .A2(G217), .A3(new_n276), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n389), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n389), .B2(new_n400), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n374), .B(new_n301), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G478), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  OAI22_X1  g225(.A1(new_n411), .A2(new_n374), .B1(KEYINPUT15), .B2(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G140), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT74), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT73), .B(G140), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G140), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT74), .B(G125), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT90), .B1(new_n424), .B2(G146), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(G125), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n415), .A2(new_n426), .A3(new_n205), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(KEYINPUT90), .A3(G146), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G237), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n276), .A3(G214), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT89), .A3(G143), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT89), .B(G143), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT18), .A2(G131), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT91), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n437), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n430), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT16), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n418), .B2(new_n423), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT16), .B1(new_n421), .B2(G125), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n445), .A2(G146), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G146), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n271), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n435), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n435), .A2(new_n453), .A3(new_n271), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT94), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(KEYINPUT94), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n443), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(new_n187), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(KEYINPUT95), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(KEYINPUT95), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n443), .B(new_n463), .C1(new_n450), .C2(new_n458), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n464), .A3(new_n301), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G475), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  INV_X1    g281(.A(new_n449), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n452), .ZN(new_n469));
  OR2_X1    g283(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n415), .A3(new_n426), .A4(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n424), .A2(KEYINPUT92), .A3(KEYINPUT19), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT92), .B1(new_n424), .B2(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n475), .B2(G146), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n461), .B1(new_n430), .B2(new_n442), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n459), .A2(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n467), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n467), .A3(new_n479), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n413), .B(new_n466), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n367), .A2(new_n373), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n314), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n487));
  INV_X1    g301(.A(new_n323), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n266), .A2(G134), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n268), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n272), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n253), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n249), .A2(new_n273), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n249), .A2(KEYINPUT66), .A3(new_n273), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT66), .B1(new_n249), .B2(new_n273), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n492), .B1(new_n227), .B2(new_n223), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n488), .B(new_n496), .C1(new_n500), .C2(KEYINPUT30), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n323), .A3(new_n495), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n431), .A2(new_n276), .A3(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n196), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT31), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n501), .A2(new_n509), .A3(new_n502), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n506), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n502), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(new_n513), .A3(new_n514), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n498), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n249), .A2(KEYINPUT66), .A3(new_n273), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n494), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n488), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n514), .B1(new_n522), .B2(new_n502), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n512), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n502), .A2(new_n513), .A3(new_n514), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n498), .A2(new_n499), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n323), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  INV_X1    g344(.A(new_n502), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT28), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT70), .A3(new_n512), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n511), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G472), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n487), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT70), .B1(new_n533), .B2(new_n512), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n525), .B(new_n506), .C1(new_n528), .C2(new_n532), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT32), .B(new_n536), .C1(new_n541), .C2(new_n511), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n323), .B1(new_n494), .B2(new_n495), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n531), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n528), .A2(new_n544), .A3(KEYINPUT29), .A4(new_n506), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n501), .A2(new_n502), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(new_n506), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n533), .A2(new_n512), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n301), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n538), .A2(new_n542), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n538), .A2(new_n542), .A3(new_n551), .A4(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n557));
  INV_X1    g371(.A(G217), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(G234), .B2(new_n301), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n203), .A2(G119), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n203), .A2(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT24), .B(G110), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT72), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n565), .B1(new_n573), .B2(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n570), .B1(new_n575), .B2(G110), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n448), .B2(new_n449), .ZN(new_n578));
  INV_X1    g392(.A(G110), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n572), .A2(new_n579), .A3(new_n574), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n569), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n427), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n449), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n564), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n576), .B1(new_n468), .B2(new_n447), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n583), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n564), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT76), .B1(new_n588), .B2(new_n564), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n587), .A2(new_n593), .A3(new_n583), .A4(new_n563), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n301), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n586), .A2(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(KEYINPUT25), .A3(new_n301), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n560), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n559), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n557), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT25), .B1(new_n599), .B2(new_n301), .ZN(new_n606));
  AND4_X1   g420(.A1(KEYINPUT25), .A2(new_n591), .A3(new_n595), .A4(new_n301), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n559), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT77), .A3(new_n603), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n486), .A2(new_n556), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND2_X1   g426(.A1(new_n605), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n535), .B2(G902), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n537), .B2(new_n535), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n309), .A2(new_n313), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n366), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n363), .B1(new_n345), .B2(new_n361), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n315), .B(new_n373), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n466), .B1(new_n482), .B2(new_n480), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n404), .B2(new_n405), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n410), .A2(new_n403), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n623), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n623), .B1(new_n410), .B2(KEYINPUT101), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n407), .A2(G902), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n411), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT102), .B(G478), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n622), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n618), .A2(new_n621), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT34), .B(G104), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n412), .A2(new_n406), .ZN(new_n644));
  INV_X1    g458(.A(new_n409), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n644), .A2(new_n645), .B1(G475), .B2(new_n465), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n478), .A2(new_n479), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n481), .A3(KEYINPUT103), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n481), .A2(KEYINPUT103), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n621), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n651), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n367), .A2(new_n653), .A3(new_n654), .A4(new_n373), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n616), .A3(new_n617), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n588), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n602), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n608), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n615), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n486), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NOR2_X1   g482(.A1(new_n372), .A2(G900), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n370), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n646), .A2(new_n649), .A3(new_n650), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n556), .A2(new_n617), .A3(new_n367), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n673), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n617), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n365), .A2(new_n366), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n547), .A2(new_n512), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n531), .A2(new_n543), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n301), .B1(new_n685), .B2(new_n506), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n538), .A2(new_n542), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n648), .A2(new_n481), .B1(G475), .B2(new_n465), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n413), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n315), .A2(new_n664), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n680), .A2(new_n681), .A3(new_n683), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  NAND3_X1  g507(.A1(new_n622), .A2(new_n639), .A3(new_n673), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n664), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n556), .A2(new_n617), .A3(new_n367), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  AOI21_X1  g511(.A(new_n613), .B1(new_n554), .B2(new_n555), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n313), .A3(new_n308), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n621), .A2(new_n640), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT41), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G113), .ZN(G15));
  NAND3_X1  g520(.A1(new_n698), .A2(new_n656), .A3(new_n702), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND2_X1  g522(.A1(new_n663), .A2(new_n484), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n701), .A2(new_n709), .A3(new_n621), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n556), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NOR2_X1   g526(.A1(new_n601), .A2(new_n604), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n528), .A2(KEYINPUT106), .A3(new_n544), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT106), .B1(new_n528), .B2(new_n544), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n506), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n536), .B1(new_n716), .B2(new_n511), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n690), .A3(new_n614), .A4(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n701), .A3(new_n621), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(G122), .Z(G24));
  NAND2_X1  g534(.A1(new_n614), .A2(new_n717), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n664), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n622), .A2(new_n639), .A3(new_n724), .A4(new_n673), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n702), .A3(new_n367), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NAND3_X1  g542(.A1(new_n365), .A2(new_n315), .A3(new_n366), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n299), .B2(G902), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n312), .B1(new_n308), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n365), .A2(new_n733), .A3(new_n315), .A4(new_n366), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT42), .B1(new_n723), .B2(new_n725), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n556), .A3(new_n610), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n726), .A2(new_n552), .A3(new_n713), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT42), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(G131), .Z(G33));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n674), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n735), .A2(new_n556), .A3(new_n610), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n283), .A2(new_n294), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n296), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n299), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n308), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT46), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n313), .B(new_n678), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n730), .A2(new_n734), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n625), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n763), .A2(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT113), .B1(new_n622), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT113), .B(KEYINPUT43), .C1(new_n622), .C2(new_n764), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n615), .A2(new_n663), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n762), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n760), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n266), .ZN(G39));
  OAI21_X1  g591(.A(new_n313), .B1(new_n756), .B2(new_n757), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(new_n313), .C1(new_n756), .C2(new_n757), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n556), .A2(new_n761), .A3(new_n610), .A4(new_n694), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  OAI211_X1 g598(.A(new_n698), .B(new_n702), .C1(new_n656), .C2(new_n703), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n719), .B1(new_n698), .B2(new_n486), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n486), .A2(new_n665), .B1(new_n710), .B2(new_n556), .ZN(new_n787));
  INV_X1    g601(.A(new_n621), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n640), .B1(new_n622), .B2(new_n413), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n616), .A2(new_n617), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n649), .A2(new_n650), .A3(new_n673), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n466), .A2(new_n792), .A3(new_n413), .A4(new_n663), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n556), .A2(new_n617), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n722), .A2(new_n726), .A3(new_n732), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n761), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n737), .A2(new_n745), .A3(new_n740), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n791), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n732), .A2(new_n367), .A3(new_n690), .ZN(new_n799));
  INV_X1    g613(.A(new_n673), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n663), .A2(KEYINPUT116), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT116), .B1(new_n663), .B2(new_n800), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(new_n801), .A3(new_n688), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n676), .A2(new_n696), .A3(new_n727), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT117), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n804), .A2(KEYINPUT117), .A3(new_n805), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT53), .B(new_n798), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n797), .A2(new_n796), .ZN(new_n812));
  INV_X1    g626(.A(new_n719), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n611), .A2(new_n666), .A3(new_n711), .A4(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n785), .A2(new_n790), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n804), .B(KEYINPUT52), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n810), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n811), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n798), .B1(new_n808), .B2(new_n809), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n819), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n779), .A2(new_n781), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n700), .A2(new_n308), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n313), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n769), .A2(new_n369), .A3(new_n368), .ZN(new_n831));
  INV_X1    g645(.A(new_n713), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n721), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n761), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n683), .A2(new_n315), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(new_n702), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT50), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n761), .A2(new_n701), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n831), .A2(new_n722), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n688), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n613), .A2(new_n370), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n844), .A2(new_n622), .A3(new_n639), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n838), .A2(KEYINPUT50), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n839), .A2(new_n841), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n825), .A2(new_n826), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n827), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n825), .B(new_n826), .C1(new_n847), .C2(new_n836), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n831), .A2(new_n367), .A3(new_n702), .A4(new_n833), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n852), .B(new_n368), .C1(new_n640), .C2(new_n844), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n831), .A2(new_n840), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n552), .A2(new_n713), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT48), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n854), .A2(KEYINPUT48), .A3(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n824), .A2(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n683), .A2(new_n622), .A3(new_n764), .A4(new_n688), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n713), .A2(new_n313), .A3(new_n315), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT114), .Z(new_n863));
  OR2_X1    g677(.A1(new_n829), .A2(KEYINPUT49), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n829), .A2(KEYINPUT49), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n276), .A2(G952), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n810), .A2(new_n818), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(G902), .ZN(new_n872));
  INV_X1    g686(.A(G210), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n336), .A2(new_n344), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n342), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT55), .Z(new_n877));
  AOI21_X1  g691(.A(new_n869), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n877), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n870), .B(new_n879), .C1(new_n872), .C2(new_n873), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(G51));
  INV_X1    g695(.A(new_n820), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n819), .B1(new_n810), .B2(new_n818), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n754), .B(KEYINPUT119), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT57), .Z(new_n886));
  OAI22_X1  g700(.A1(new_n884), .A2(new_n886), .B1(new_n307), .B2(new_n306), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n753), .B(KEYINPUT120), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n871), .A2(G902), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n869), .B1(new_n887), .B2(new_n891), .ZN(G54));
  NAND2_X1  g706(.A1(KEYINPUT58), .A2(G475), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n301), .B(new_n893), .C1(new_n810), .C2(new_n818), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT122), .B1(new_n894), .B2(new_n478), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n869), .B1(new_n894), .B2(new_n478), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n894), .A2(KEYINPUT122), .A3(new_n478), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(G60));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n763), .B1(new_n824), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n869), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n763), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n884), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(G63));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n910));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n871), .A2(new_n661), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n904), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n810), .B2(new_n818), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n599), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n909), .B(new_n910), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n916), .A2(new_n599), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n869), .B1(new_n916), .B2(new_n661), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT123), .A4(new_n908), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n918), .A2(new_n921), .ZN(G66));
  INV_X1    g736(.A(new_n371), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n923), .B2(new_n339), .ZN(new_n924));
  INV_X1    g738(.A(new_n791), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n875), .B1(G898), .B2(new_n276), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT124), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  OR2_X1    g743(.A1(new_n500), .A2(KEYINPUT30), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n496), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n475), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT127), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n932), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n797), .B(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n367), .A2(new_n690), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n774), .B1(new_n855), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n760), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n676), .A2(new_n727), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n783), .A2(new_n696), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n276), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n276), .A2(G900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT126), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n937), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n692), .A2(new_n696), .A3(new_n942), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n698), .A2(new_n762), .A3(new_n789), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n783), .B1(new_n679), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n776), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n932), .B1(new_n957), .B2(new_n276), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n936), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(new_n950), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n949), .B1(new_n945), .B2(new_n946), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n932), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n963), .A3(new_n935), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n957), .B2(new_n791), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n869), .B1(new_n968), .B2(new_n684), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n547), .A2(new_n506), .ZN(new_n970));
  INV_X1    g784(.A(new_n507), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n823), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n967), .B1(new_n944), .B2(new_n791), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n547), .A3(new_n512), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n969), .A2(new_n973), .A3(new_n975), .ZN(G57));
endmodule


