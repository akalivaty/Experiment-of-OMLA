//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n536,
    new_n537, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  OAI21_X1  g032(.A(KEYINPUT67), .B1(new_n457), .B2(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n457), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n462));
  NAND4_X1  g037(.A1(new_n460), .A2(G137), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n457), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n459), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n459), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n474), .B2(G2105), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n460), .A2(G2105), .A3(new_n462), .ZN(new_n481));
  OAI221_X1 g056(.A(new_n477), .B1(new_n478), .B2(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n460), .A2(G126), .A3(G2105), .A4(new_n462), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n460), .A2(G138), .A3(new_n461), .A4(new_n462), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n470), .B2(new_n471), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n489), .B2(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT5), .B(G543), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G88), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G50), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n494), .A2(G62), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(KEYINPUT68), .B1(G75), .B2(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(KEYINPUT68), .B2(new_n501), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n500), .B1(new_n503), .B2(G651), .ZN(G166));
  AND2_X1   g079(.A1(G63), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n506));
  NAND3_X1  g081(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n494), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n495), .A2(G51), .A3(G543), .ZN(new_n511));
  INV_X1    g086(.A(G89), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n496), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n510), .A2(new_n513), .ZN(G168));
  NAND3_X1  g089(.A1(new_n495), .A2(G52), .A3(G543), .ZN(new_n515));
  INV_X1    g090(.A(G90), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n496), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n522), .A3(G64), .ZN(new_n523));
  NAND2_X1  g098(.A1(G77), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n525), .ZN(G171));
  AOI22_X1  g101(.A1(new_n494), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n518), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n495), .A2(G43), .A3(G543), .ZN(new_n529));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n496), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G860), .ZN(G153));
  AND3_X1   g108(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G36), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT8), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G188));
  AND2_X1   g113(.A1(new_n495), .A2(G543), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT69), .B(KEYINPUT9), .Z(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G53), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n542));
  INV_X1    g117(.A(G53), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n498), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n494), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G91), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n546), .A2(new_n518), .B1(new_n496), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n545), .A2(new_n548), .ZN(G299));
  INV_X1    g124(.A(G171), .ZN(G301));
  NAND2_X1  g125(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  AND4_X1   g128(.A1(new_n520), .A2(new_n522), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G89), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n555), .A2(new_n509), .A3(new_n508), .A4(new_n511), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  OAI21_X1  g132(.A(G651), .B1(new_n494), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n554), .A2(G87), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n495), .A2(G49), .A3(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT70), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n494), .B2(G61), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n565), .B1(new_n568), .B2(new_n518), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n520), .A2(new_n522), .A3(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(new_n566), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT72), .A3(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n554), .A2(G86), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n551), .A2(new_n553), .A3(G48), .A4(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n495), .A2(KEYINPUT73), .A3(G48), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n569), .A2(new_n572), .A3(new_n573), .A4(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n539), .A2(G47), .B1(new_n554), .B2(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n494), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n518), .B2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n496), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n554), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n520), .A2(new_n522), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(G651), .A2(new_n592), .B1(new_n539), .B2(G54), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n583), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n583), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n545), .A2(new_n548), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT74), .Z(G297));
  XOR2_X1   g175(.A(new_n599), .B(KEYINPUT75), .Z(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n594), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n594), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n532), .ZN(new_n606));
  MUX2_X1   g181(.A(new_n605), .B(new_n606), .S(KEYINPUT76), .Z(G323));
  XNOR2_X1  g182(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n608));
  XNOR2_X1  g183(.A(G323), .B(new_n608), .ZN(G282));
  INV_X1    g184(.A(new_n481), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G123), .ZN(new_n611));
  INV_X1    g186(.A(new_n478), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n461), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NOR2_X1   g192(.A1(new_n467), .A2(G2104), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT66), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n459), .A2(new_n468), .A3(new_n469), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n464), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT13), .B(G2100), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n617), .A2(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(KEYINPUT80), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n629), .A2(new_n630), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT81), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n657), .A2(KEYINPUT17), .A3(new_n654), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n657), .B2(KEYINPUT17), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n658), .A2(new_n659), .A3(new_n653), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR3_X1    g247(.A1(new_n669), .A2(KEYINPUT82), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(KEYINPUT82), .B1(new_n669), .B2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT20), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  MUX2_X1   g252(.A(new_n676), .B(new_n677), .S(new_n669), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(KEYINPUT20), .B1(new_n673), .B2(new_n674), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n679), .A2(G1991), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(G1991), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  AOI21_X1  g257(.A(G1996), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(G1996), .A3(new_n682), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n667), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n685), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n687), .A2(new_n666), .A3(new_n683), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n665), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n666), .B1(new_n687), .B2(new_n683), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n667), .A3(new_n685), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n691), .A3(new_n664), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G6), .ZN(new_n704));
  INV_X1    g279(.A(G305), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n698), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT34), .Z(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(G1986), .Z(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT83), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n610), .A2(G119), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n612), .A2(G131), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n710), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n699), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n699), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT87), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1966), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT88), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT31), .B(G11), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT89), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G28), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n713), .B1(new_n734), .B2(G28), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n735), .B2(new_n736), .C1(new_n616), .C2(new_n713), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT90), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n729), .A2(G1966), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G171), .B2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n739), .B1(G1961), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n731), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT91), .Z(new_n744));
  INV_X1    g319(.A(KEYINPUT23), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n745), .A2(new_n699), .A3(G20), .ZN(new_n746));
  NAND2_X1  g321(.A1(G299), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n745), .B1(new_n699), .B2(G20), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n713), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n713), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT29), .B(G2090), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n464), .A2(G103), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n622), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n759), .B1(new_n760), .B2(new_n478), .C1(new_n761), .C2(new_n461), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(G29), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n612), .A2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n610), .A2(G129), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n770), .A2(new_n771), .B1(G105), .B2(new_n464), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n766), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G29), .B2(G32), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n713), .B1(KEYINPUT24), .B2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(KEYINPUT24), .B2(G34), .ZN(new_n780));
  INV_X1    g355(.A(G160), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n764), .A2(G2072), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n765), .A2(new_n778), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n776), .A2(new_n777), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n699), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n594), .B2(new_n699), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n699), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n532), .B2(new_n699), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT84), .B(G1341), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n793), .A2(new_n795), .B1(new_n741), .B2(G1961), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n782), .A2(new_n783), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n787), .A2(new_n791), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n713), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n713), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n756), .A2(new_n786), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n713), .A2(G26), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n610), .A2(KEYINPUT85), .A3(G128), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n612), .A2(G140), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT85), .ZN(new_n808));
  INV_X1    g383(.A(G128), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n481), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n806), .A2(new_n807), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n804), .B(new_n805), .C1(new_n813), .C2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n804), .B2(new_n805), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT86), .B(G2067), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n726), .A2(new_n744), .A3(new_n818), .ZN(G311));
  NOR2_X1   g394(.A1(new_n744), .A2(new_n818), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n724), .B(KEYINPUT36), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n590), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G651), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n554), .A2(G93), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT93), .B(G55), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n495), .A2(new_n828), .A3(G543), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n594), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT95), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n829), .B1(new_n496), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n494), .A2(G67), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n518), .B1(new_n839), .B2(new_n823), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT94), .A4(new_n829), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n532), .A3(new_n842), .ZN(new_n843));
  OAI221_X1 g418(.A(new_n529), .B1(new_n496), .B2(new_n530), .C1(new_n527), .C2(new_n518), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(new_n830), .A3(new_n836), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n835), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT96), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n833), .B1(new_n852), .B2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(new_n781), .B(new_n616), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n610), .A2(G130), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n612), .A2(G142), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n720), .A2(new_n864), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n867), .A2(new_n868), .A3(new_n625), .ZN(new_n869));
  INV_X1    g444(.A(new_n625), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n720), .A2(new_n864), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n625), .B1(new_n867), .B2(new_n868), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n871), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(KEYINPUT99), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n489), .A2(new_n492), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n484), .A2(KEYINPUT98), .A3(new_n486), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT98), .B1(new_n484), .B2(new_n486), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(new_n813), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n813), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n773), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n773), .A3(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n763), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n762), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n878), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n878), .B1(new_n890), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n890), .B(new_n888), .C1(new_n869), .C2(new_n873), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n890), .A2(new_n888), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n895), .B(new_n857), .C1(new_n896), .C2(new_n878), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT40), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(G395));
  NAND2_X1  g482(.A1(G299), .A2(new_n594), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n588), .A2(new_n593), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n598), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n604), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n846), .ZN(new_n918));
  MUX2_X1   g493(.A(new_n915), .B(new_n911), .S(new_n918), .Z(new_n919));
  XNOR2_X1  g494(.A(G166), .B(G288), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n705), .B(G290), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n920), .B(new_n921), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n926), .A2(KEYINPUT103), .B1(KEYINPUT42), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n919), .A2(KEYINPUT104), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n927), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n931), .B2(new_n919), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT104), .B1(new_n931), .B2(new_n919), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G868), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n830), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n517), .B2(new_n525), .ZN(new_n942));
  INV_X1    g517(.A(new_n525), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n554), .A2(G90), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT105), .A4(new_n515), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n945), .A3(G286), .ZN(new_n946));
  NAND3_X1  g521(.A1(G168), .A2(G171), .A3(KEYINPUT105), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n843), .A2(new_n946), .A3(new_n947), .A4(new_n845), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n845), .A2(new_n843), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT106), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n949), .A2(new_n950), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n954), .A2(new_n915), .B1(new_n911), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n928), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n946), .A2(new_n947), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n846), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n952), .B1(new_n959), .B2(new_n948), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n948), .A2(new_n952), .ZN(new_n961));
  INV_X1    g536(.A(new_n911), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n913), .A2(new_n914), .B1(new_n959), .B2(new_n948), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n924), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT107), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n924), .B(new_n967), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n957), .A2(new_n966), .A3(KEYINPUT43), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n915), .B1(new_n960), .B2(new_n961), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n955), .A2(new_n911), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n928), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n894), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n928), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n940), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n957), .A2(new_n966), .A3(new_n970), .A4(new_n968), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n940), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n939), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT44), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n977), .A2(new_n984), .A3(KEYINPUT108), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(G397));
  XNOR2_X1  g561(.A(KEYINPUT109), .B(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n882), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  INV_X1    g564(.A(G125), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n620), .B2(new_n621), .ZN(new_n991));
  INV_X1    g566(.A(new_n473), .ZN(new_n992));
  OAI21_X1  g567(.A(G2105), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n466), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n993), .A2(G40), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT111), .B1(new_n999), .B2(G1996), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n997), .A2(new_n1001), .A3(new_n1002), .A4(new_n998), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n773), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n813), .B(G2067), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n773), .A2(G1996), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n999), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n720), .B(new_n722), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n695), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT116), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n569), .A2(new_n1018), .A3(new_n572), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G1981), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT72), .B1(new_n571), .B2(G651), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n565), .B(new_n518), .C1(new_n570), .C2(new_n566), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n576), .A2(new_n577), .B1(new_n554), .B2(G86), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND4_X1   g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n572), .A4(new_n569), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1020), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n882), .A2(G40), .A3(new_n1029), .A4(G160), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n1024), .B2(new_n1018), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1028), .A2(G8), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1017), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n705), .A2(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT117), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(G8), .A3(new_n1030), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n560), .A2(new_n563), .A3(G1976), .A4(new_n561), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1030), .A2(G8), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(new_n1030), .A3(G8), .A4(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1046), .A3(new_n1036), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1044), .A2(new_n1036), .A3(new_n1049), .A4(new_n1046), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G166), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT113), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1057), .A3(KEYINPUT55), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n993), .A2(G40), .A3(new_n994), .ZN(new_n1060));
  AOI22_X1  g635(.A1(KEYINPUT4), .A2(new_n488), .B1(new_n622), .B2(new_n491), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1029), .B1(new_n1061), .B2(new_n487), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(KEYINPUT50), .ZN(new_n1063));
  INV_X1    g638(.A(G2090), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n882), .A2(new_n1065), .A3(new_n1029), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1060), .B1(new_n1062), .B2(new_n989), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1971), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT112), .B(G1971), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1059), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1040), .A2(new_n1041), .B1(new_n1051), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1055), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n995), .B1(new_n1062), .B2(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1065), .B1(new_n882), .B2(new_n1029), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1077), .A2(new_n1078), .A3(G2090), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1047), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1063), .A2(new_n1083), .A3(new_n1066), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n995), .B1(new_n1062), .B2(new_n989), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT45), .B1(new_n882), .B2(new_n1029), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(G2078), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n989), .B1(G164), .B2(G1384), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1069), .A2(new_n1092), .A3(new_n1093), .A4(new_n995), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1089), .A2(new_n1091), .B1(new_n1094), .B2(new_n1090), .ZN(new_n1095));
  AOI21_X1  g670(.A(G301), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1081), .A2(new_n1074), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1063), .A2(new_n783), .A3(new_n1066), .ZN(new_n1098));
  OAI211_X1 g673(.A(G168), .B(new_n1098), .C1(new_n1089), .C2(G1966), .ZN(new_n1099));
  AND2_X1   g674(.A1(KEYINPUT124), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1098), .B1(new_n1089), .B2(G1966), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(G8), .A3(G286), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(new_n1105), .A3(new_n1100), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1097), .B1(KEYINPUT62), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(new_n1109), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1075), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1069), .ZN(new_n1113));
  INV_X1    g688(.A(new_n487), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1384), .B1(new_n879), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n995), .B1(new_n1115), .B2(KEYINPUT45), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n702), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1067), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1059), .B1(new_n1120), .B2(G8), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1112), .B1(new_n1121), .B2(new_n1051), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1076), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT118), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1103), .A2(G8), .A3(G168), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(new_n1074), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1122), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1081), .A2(new_n1074), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1131), .B2(new_n1126), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(G171), .B(KEYINPUT54), .Z(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1086), .A2(KEYINPUT125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1094), .A2(new_n1090), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n988), .A2(new_n989), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n995), .A3(new_n1091), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1139), .B(new_n1136), .C1(new_n1113), .C2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1086), .A2(KEYINPUT125), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1137), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1131), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1107), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1030), .A2(G2067), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT121), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1063), .A2(new_n1083), .A3(new_n1066), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1152), .B2(new_n790), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n909), .B1(new_n1153), .B2(KEYINPUT60), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1348), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NOR4_X1   g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n594), .A4(new_n1148), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1154), .A2(new_n1157), .B1(KEYINPUT60), .B2(new_n1153), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n750), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT119), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT120), .Z(new_n1162));
  OR2_X1    g737(.A1(new_n1160), .A2(KEYINPUT119), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(G299), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1163), .B(new_n1162), .C1(new_n545), .C2(new_n548), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1068), .A2(new_n1069), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1159), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1159), .B2(new_n1169), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1176), .B(new_n1172), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1173), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(G1996), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1068), .A2(KEYINPUT122), .A3(new_n1002), .A4(new_n1069), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT58), .B(G1341), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n1030), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n532), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1188), .A3(new_n532), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1158), .A2(new_n1178), .A3(new_n1190), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1153), .A2(new_n909), .A3(new_n1170), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1192), .A2(new_n1171), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1147), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1014), .B1(new_n1134), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n720), .A2(new_n722), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT126), .Z(new_n1197));
  NOR3_X1   g772(.A1(new_n1004), .A2(new_n1007), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n813), .A2(G2067), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1009), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n999), .A2(G1986), .A3(G290), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT48), .Z(new_n1202));
  NAND3_X1  g777(.A1(new_n1202), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT46), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1000), .A2(KEYINPUT46), .A3(new_n1003), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1005), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1009), .B1(new_n773), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1204), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1000), .A2(KEYINPUT46), .A3(new_n1003), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT46), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n1204), .B(new_n1211), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1215), .ZN(new_n1216));
  OAI211_X1 g791(.A(new_n1200), .B(new_n1203), .C1(new_n1212), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1195), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g794(.A(G319), .ZN(new_n1221));
  AOI211_X1 g795(.A(new_n1221), .B(G227), .C1(new_n647), .C2(new_n649), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n689), .A2(new_n1222), .A3(new_n692), .ZN(new_n1223));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g799(.A1(new_n689), .A2(new_n1222), .A3(KEYINPUT127), .A4(new_n692), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n1225), .A2(new_n981), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n905), .B2(new_n903), .ZN(G308));
  XNOR2_X1  g802(.A(new_n898), .B(new_n899), .ZN(new_n1229));
  NAND4_X1  g803(.A1(new_n1229), .A2(new_n981), .A3(new_n1225), .A4(new_n1226), .ZN(G225));
endmodule


