//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  OR3_X1    g0017(.A1(new_n206), .A2(KEYINPUT65), .A3(G13), .ZN(new_n218));
  OAI21_X1  g0018(.A(KEYINPUT65), .B1(new_n206), .B2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT0), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n217), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1698), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n248), .B2(new_n249), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n255), .A2(G223), .B1(new_n258), .B2(G77), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n247), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n247), .A3(G274), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n247), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n264), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G190), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n225), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n226), .B1(new_n201), .B2(new_n203), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n226), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n226), .A2(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n273), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n273), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n226), .B2(G1), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n266), .A2(KEYINPUT68), .A3(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n284), .A2(G50), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n281), .B(new_n289), .C1(G50), .C2(new_n282), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n271), .B(new_n291), .C1(new_n292), .C2(new_n270), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n270), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n260), .B2(new_n269), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n265), .A2(new_n254), .ZN(new_n303));
  INV_X1    g0103(.A(G232), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G1698), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n305), .C1(new_n256), .C2(new_n257), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n247), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n247), .A2(G238), .A3(new_n267), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n264), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(KEYINPUT13), .C1(new_n308), .C2(new_n311), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT13), .B1(new_n308), .B2(new_n311), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n317), .A2(KEYINPUT72), .A3(G179), .A4(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(G179), .A3(new_n314), .A4(new_n316), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n299), .B1(new_n314), .B2(new_n318), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT14), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n226), .A2(G33), .A3(G77), .ZN(new_n328));
  INV_X1    g0128(.A(G50), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n328), .B1(new_n226), .B2(G68), .C1(new_n279), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n273), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT11), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n282), .A2(G68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n284), .A2(G68), .A3(new_n288), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n334), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n314), .A2(new_n318), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n341), .B2(G200), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n319), .A2(G190), .A3(new_n314), .A4(new_n316), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n342), .A2(KEYINPUT71), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT71), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G244), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n264), .B1(new_n348), .B2(new_n268), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n250), .A2(G232), .B1(new_n258), .B2(G107), .ZN(new_n350));
  INV_X1    g0150(.A(new_n255), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n209), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n247), .B1(new_n352), .B2(KEYINPUT69), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n350), .B(new_n354), .C1(new_n209), .C2(new_n351), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n288), .A2(G77), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n284), .B1(new_n202), .B2(new_n283), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n275), .A2(new_n279), .B1(new_n226), .B2(new_n202), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n276), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n273), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n356), .B2(G169), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(G200), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n366), .B1(new_n356), .B2(G190), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT3), .B(G33), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n208), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n208), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n203), .ZN(new_n380));
  INV_X1    g0180(.A(new_n279), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n372), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n258), .B2(new_n226), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n256), .A2(new_n257), .A3(new_n373), .A4(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n383), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n389), .A3(new_n273), .ZN(new_n390));
  INV_X1    g0190(.A(new_n275), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n284), .A2(new_n288), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n283), .B2(new_n275), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n278), .A2(new_n210), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G223), .A2(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n265), .B2(G1698), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(new_n374), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT73), .B1(new_n398), .B2(new_n247), .ZN(new_n399));
  OR2_X1    g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n265), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n256), .C2(new_n257), .ZN(new_n402));
  INV_X1    g0202(.A(new_n395), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n247), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n247), .A2(G232), .A3(new_n267), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n264), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n299), .B1(new_n404), .B2(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n394), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT18), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n390), .B2(new_n393), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n408), .A2(G190), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n399), .A2(new_n406), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n292), .B1(new_n404), .B2(new_n408), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n390), .A2(new_n423), .A3(new_n393), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n390), .A2(new_n423), .A3(new_n393), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n371), .A2(new_n419), .A3(new_n429), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n302), .A2(new_n347), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT84), .ZN(new_n432));
  INV_X1    g0232(.A(new_n247), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n266), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(KEYINPUT76), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(KEYINPUT76), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT83), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n374), .A2(KEYINPUT83), .A3(G257), .A4(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G294), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n374), .A2(G250), .A3(new_n254), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n439), .A2(G264), .B1(new_n446), .B2(new_n433), .ZN(new_n447));
  INV_X1    g0247(.A(G274), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n433), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n437), .A2(new_n449), .A3(new_n438), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n299), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n433), .ZN(new_n452));
  INV_X1    g0252(.A(new_n438), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(new_n247), .C1(new_n453), .C2(new_n436), .ZN(new_n454));
  AND4_X1   g0254(.A1(G179), .A2(new_n452), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n432), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n450), .A3(new_n454), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G169), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(KEYINPUT84), .C1(new_n297), .C2(new_n457), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n226), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n374), .A2(new_n462), .A3(new_n226), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n278), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n226), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n226), .B2(G107), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(KEYINPUT23), .A3(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n464), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n473), .A2(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n467), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n461), .B2(new_n463), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT24), .B1(new_n479), .B2(KEYINPUT81), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n476), .B(new_n273), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n272), .A2(new_n225), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n266), .A2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n282), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n470), .B1(KEYINPUT82), .B2(KEYINPUT25), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n282), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n283), .A2(KEYINPUT82), .A3(KEYINPUT25), .A4(new_n470), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n485), .A2(G107), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n456), .A2(new_n459), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT85), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n484), .A2(new_n363), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n363), .A2(new_n283), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT19), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n226), .B1(new_n307), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n210), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n226), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n500), .B1(new_n276), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT77), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n482), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT77), .A4(new_n507), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n497), .B(new_n499), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n211), .B1(new_n262), .B2(G1), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n266), .A2(new_n448), .A3(G45), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n247), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n516));
  OAI211_X1 g0316(.A(G238), .B(new_n254), .C1(new_n256), .C2(new_n257), .ZN(new_n517));
  INV_X1    g0317(.A(new_n466), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(new_n433), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n297), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G169), .B2(new_n520), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n433), .ZN(new_n523));
  INV_X1    g0323(.A(new_n515), .ZN(new_n524));
  AOI21_X1  g0324(.A(G200), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(G190), .B(new_n515), .C1(new_n519), .C2(new_n433), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n508), .A2(new_n509), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n273), .A3(new_n511), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n485), .A2(G87), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n498), .A3(new_n530), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n512), .A2(new_n522), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n481), .A2(new_n490), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n457), .A2(new_n292), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G190), .B2(new_n457), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT21), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT78), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n255), .A2(new_n538), .A3(G264), .ZN(new_n539));
  OAI211_X1 g0339(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n250), .A2(G257), .B1(new_n258), .B2(G303), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n247), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G270), .B(new_n247), .C1(new_n453), .C2(new_n436), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n450), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G169), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT79), .B1(new_n484), .B2(new_n465), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n284), .A2(new_n549), .A3(G116), .A4(new_n483), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n282), .A2(G116), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n226), .C1(G33), .C2(new_n506), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n465), .A2(G20), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n273), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT20), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n537), .B1(new_n547), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n542), .A2(new_n543), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n433), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n450), .A2(new_n545), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(G190), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n544), .B2(new_n546), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n563), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n551), .B(new_n554), .C1(new_n560), .C2(new_n561), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT21), .A4(G169), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n544), .A2(new_n546), .A3(new_n297), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n572), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n564), .A2(new_n570), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n282), .A2(G97), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n485), .B2(G97), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G107), .B1(new_n385), .B2(new_n386), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g0383(.A(KEYINPUT74), .B(G107), .Z(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g0385(.A(KEYINPUT74), .B(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n582), .A3(new_n581), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(G20), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n381), .A2(G77), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n579), .B1(new_n590), .B2(new_n273), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(new_n247), .C1(new_n453), .C2(new_n436), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n450), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(new_n254), .C1(new_n256), .C2(new_n257), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n374), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n374), .A2(G250), .A3(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n555), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n433), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(G190), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n591), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n599), .A2(KEYINPUT75), .A3(new_n433), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT75), .B1(new_n599), .B2(new_n433), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n593), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n593), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n590), .A2(new_n273), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n299), .B1(new_n608), .B2(new_n578), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n297), .B(new_n593), .C1(new_n603), .C2(new_n604), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n602), .A2(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n536), .A2(new_n576), .A3(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n431), .A2(new_n496), .A3(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n301), .ZN(new_n614));
  INV_X1    g0414(.A(new_n368), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n344), .A2(new_n345), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n340), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n429), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n419), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n614), .B1(new_n619), .B2(new_n296), .ZN(new_n620));
  AOI21_X1  g0420(.A(G200), .B1(new_n447), .B2(new_n450), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n457), .A2(G190), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n481), .B(new_n490), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n450), .A2(new_n592), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT75), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n600), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n599), .A2(KEYINPUT75), .A3(new_n433), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n591), .B(new_n601), .C1(new_n628), .C2(new_n292), .ZN(new_n629));
  INV_X1    g0429(.A(new_n600), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n299), .B1(new_n630), .B2(new_n624), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n608), .A2(new_n578), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n610), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n529), .A2(new_n498), .A3(new_n530), .ZN(new_n634));
  INV_X1    g0434(.A(G190), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n520), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(G200), .B2(new_n520), .ZN(new_n637));
  AOI21_X1  g0437(.A(G169), .B1(new_n523), .B2(new_n524), .ZN(new_n638));
  AOI211_X1 g0438(.A(G179), .B(new_n515), .C1(new_n519), .C2(new_n433), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n497), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n529), .A2(new_n641), .A3(new_n498), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n634), .A2(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n623), .A2(new_n629), .A3(new_n633), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n564), .A2(new_n573), .A3(new_n575), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n458), .B1(new_n297), .B2(new_n457), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n491), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n633), .B2(new_n532), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n643), .A2(new_n651), .A3(new_n610), .A4(new_n609), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n512), .A2(new_n522), .ZN(new_n655));
  INV_X1    g0455(.A(new_n633), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n643), .ZN(new_n657));
  NOR2_X1   g0457(.A1(KEYINPUT86), .A2(KEYINPUT26), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n654), .A2(KEYINPUT87), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n650), .B2(new_n652), .ZN(new_n663));
  INV_X1    g0463(.A(new_n655), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n633), .A2(new_n532), .ZN(new_n665));
  INV_X1    g0465(.A(new_n658), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n661), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n649), .B1(new_n660), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n620), .B1(new_n431), .B2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n266), .A2(new_n226), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT88), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n481), .B2(new_n490), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n533), .B2(new_n535), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n494), .A2(new_n495), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n492), .A2(new_n676), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n679), .A2(KEYINPUT90), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT90), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n676), .A2(new_n563), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n645), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT89), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n564), .A2(new_n570), .A3(new_n573), .A4(new_n575), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n685), .B(KEYINPUT89), .C1(new_n687), .C2(new_n684), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n688), .A3(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n676), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n646), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n679), .A2(new_n680), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n679), .A2(KEYINPUT90), .A3(new_n680), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n648), .A2(new_n692), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n691), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n220), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n502), .A2(new_n210), .A3(new_n465), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n704), .A2(new_n266), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n224), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NOR3_X1   g0508(.A1(new_n669), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n494), .A2(new_n495), .A3(new_n646), .ZN(new_n710));
  INV_X1    g0510(.A(new_n644), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n653), .A2(new_n655), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n692), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n644), .A2(new_n687), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n494), .A3(new_n495), .A4(new_n676), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n447), .A2(new_n593), .A3(new_n600), .A4(new_n520), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n566), .A2(new_n567), .A3(G179), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n593), .A2(new_n600), .A3(new_n520), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n574), .A3(KEYINPUT30), .A4(new_n447), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n520), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n605), .A2(new_n457), .A3(new_n571), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n728), .B2(new_n692), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n717), .B1(new_n719), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n709), .A2(new_n716), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n708), .B1(new_n733), .B2(G1), .ZN(G364));
  AND2_X1   g0534(.A1(new_n226), .A2(G13), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n266), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n704), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n689), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(G330), .B1(new_n686), .B2(new_n688), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n686), .B2(new_n688), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n703), .A2(new_n374), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n224), .A2(new_n262), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(new_n262), .C2(new_n244), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n220), .A2(G355), .A3(new_n374), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n750), .C1(G116), .C2(new_n220), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n225), .B1(G20), .B2(new_n299), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n739), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n635), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n226), .A2(new_n635), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n297), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n759), .A2(new_n329), .B1(new_n762), .B2(new_n378), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n226), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n761), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n763), .B1(new_n771), .B2(G77), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n292), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n760), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G87), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n764), .A2(new_n779), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n374), .C1(new_n470), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n226), .B1(new_n774), .B2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n757), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n789), .B2(new_n208), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n778), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n258), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n759), .A2(new_n794), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n793), .B(new_n796), .C1(new_n788), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n776), .A2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n780), .C1(new_n801), .C2(new_n762), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G311), .B2(new_n771), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n773), .A2(new_n791), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n752), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n756), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n740), .A2(new_n741), .B1(new_n746), .B2(new_n806), .ZN(G396));
  INV_X1    g0607(.A(new_n762), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G143), .B1(G137), .B2(new_n758), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n277), .B2(new_n789), .C1(new_n770), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  NOR2_X1   g0612(.A1(new_n785), .A2(new_n378), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n374), .B1(new_n780), .B2(new_n329), .ZN(new_n814));
  INV_X1    g0614(.A(new_n783), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G68), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n775), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n770), .A2(new_n465), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT94), .B(G283), .Z(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n822), .A2(new_n788), .B1(new_n758), .B2(G303), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n374), .B1(new_n776), .B2(G311), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n787), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n783), .A2(new_n210), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n470), .A2(new_n780), .B1(new_n762), .B2(new_n795), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n820), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n752), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n752), .A2(new_n742), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n739), .B1(new_n202), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n358), .A2(new_n367), .A3(new_n692), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n369), .A2(new_n370), .ZN(new_n833));
  INV_X1    g0633(.A(new_n366), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n676), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(new_n835), .B2(new_n615), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n829), .B(new_n831), .C1(new_n836), .C2(new_n743), .ZN(new_n837));
  INV_X1    g0637(.A(new_n649), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT87), .B1(new_n654), .B2(new_n659), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n663), .A2(new_n667), .A3(new_n661), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n836), .B1(new_n841), .B2(new_n676), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT95), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n371), .A2(new_n676), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n669), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(KEYINPUT95), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n732), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n739), .B1(new_n848), .B2(new_n732), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n837), .B1(new_n850), .B2(new_n851), .ZN(G384));
  NAND2_X1  g0652(.A1(new_n585), .A2(new_n587), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  OAI211_X1 g0654(.A(G116), .B(new_n227), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n201), .A2(G68), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(KEYINPUT96), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n379), .A2(new_n223), .A3(new_n202), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n858), .B2(KEYINPUT96), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n266), .B(G13), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n302), .A2(new_n430), .A3(new_n347), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n709), .B2(new_n716), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n620), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT102), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n832), .A2(KEYINPUT97), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n832), .A2(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT98), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT98), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT95), .B1(new_n841), .B2(new_n846), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n669), .A2(new_n843), .A3(new_n844), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n415), .A2(new_n425), .A3(new_n418), .A4(new_n428), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n394), .A3(new_n675), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n394), .A2(new_n675), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n414), .A2(new_n881), .A3(new_n426), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n414), .A2(new_n881), .A3(new_n884), .A4(new_n426), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n880), .B2(new_n886), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n339), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n676), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n347), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n340), .A2(new_n346), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n878), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n419), .A2(new_n675), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n887), .A2(new_n888), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n424), .A2(new_n416), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n903), .A2(KEYINPUT100), .A3(new_n884), .A4(new_n881), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n904), .A3(new_n883), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT101), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n902), .A2(new_n904), .A3(new_n883), .A4(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n880), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n900), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n887), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n899), .B1(new_n912), .B2(new_n898), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n890), .B1(new_n324), .B2(new_n326), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n676), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT99), .Z(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n897), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n896), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n867), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n719), .A2(new_n731), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n836), .A3(new_n895), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n887), .B2(new_n888), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n893), .B1(new_n340), .B2(new_n346), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n914), .A2(new_n616), .A3(new_n891), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n836), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n719), .B2(new_n731), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n908), .A2(new_n880), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n905), .A2(new_n906), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n932), .B2(new_n887), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n933), .B2(KEYINPUT40), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n864), .A2(new_n921), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n717), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n266), .B2(new_n735), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n920), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n863), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI21_X1  g0742(.A(new_n755), .B1(new_n220), .B2(new_n363), .ZN(new_n943));
  INV_X1    g0743(.A(new_n747), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n237), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n738), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT110), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n771), .A2(new_n822), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n780), .A2(new_n465), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(KEYINPUT46), .B1(new_n470), .B2(new_n785), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G311), .B2(new_n758), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n783), .A2(new_n506), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n258), .B1(new_n762), .B2(new_n800), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G317), .C2(new_n776), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n949), .A2(KEYINPUT46), .B1(G294), .B2(new_n788), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n948), .A2(new_n951), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n201), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n771), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n374), .B1(new_n762), .B2(new_n277), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G159), .B2(new_n788), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n786), .A2(G68), .B1(G143), .B2(new_n758), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n783), .A2(new_n202), .B1(new_n775), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G58), .B2(new_n781), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n965), .A3(KEYINPUT47), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT47), .B1(new_n956), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n805), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n947), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n692), .A2(new_n531), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n643), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n664), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n969), .B1(new_n745), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n632), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n629), .A2(new_n974), .A3(new_n633), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT104), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n611), .A2(KEYINPUT104), .A3(new_n974), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n633), .C2(new_n676), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n690), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT108), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n693), .B(new_n979), .C1(new_n681), .C2(new_n682), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n977), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n656), .B1(new_n985), .B2(new_n496), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n692), .B1(new_n986), .B2(KEYINPUT105), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n983), .A2(KEYINPUT42), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n984), .B1(new_n989), .B2(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT106), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n972), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n990), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n990), .A2(new_n994), .A3(KEYINPUT107), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n997), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n990), .B2(new_n994), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n982), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n981), .B(new_n1005), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n693), .B1(new_n681), .B2(new_n682), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n700), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n979), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n979), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1019), .B(new_n979), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1014), .A2(new_n1015), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n690), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n683), .A2(new_n694), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n689), .B(KEYINPUT109), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1023), .A2(new_n1024), .A3(new_n1010), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n689), .A2(KEYINPUT109), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1023), .B2(new_n1010), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(new_n733), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n701), .B2(new_n979), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1016), .A2(KEYINPUT44), .A3(new_n1017), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1012), .B(new_n1013), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n691), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1022), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n733), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n704), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n737), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n973), .B1(new_n1009), .B2(new_n1039), .ZN(G387));
  INV_X1    g0840(.A(new_n704), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1029), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n733), .B2(new_n1028), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1028), .A2(new_n737), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n258), .B1(new_n775), .B2(new_n794), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n808), .A2(G317), .B1(G311), .B2(new_n788), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n801), .B2(new_n759), .C1(new_n770), .C2(new_n800), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n786), .A2(new_n822), .B1(new_n781), .B2(G294), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  AOI211_X1 g0853(.A(new_n1045), .B(new_n1053), .C1(G116), .C2(new_n815), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n781), .A2(G77), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n277), .B2(new_n775), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1056), .A2(new_n258), .A3(new_n952), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT111), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n785), .A2(new_n363), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n808), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n391), .A2(new_n788), .B1(G159), .B2(new_n758), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n770), .C2(new_n208), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n752), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n683), .A2(new_n744), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n234), .A2(new_n262), .A3(new_n374), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n275), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n275), .B2(G50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n705), .B1(new_n1070), .B2(new_n258), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n220), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n754), .B1(G107), .B2(new_n703), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n739), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1064), .A2(new_n1065), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1043), .A2(new_n1044), .A3(new_n1075), .ZN(G393));
  INV_X1    g0876(.A(new_n1029), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1021), .A2(new_n690), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n691), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n704), .A3(new_n1035), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n755), .B1(new_n506), .B2(new_n220), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n944), .A2(new_n241), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n738), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n979), .A2(new_n745), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n759), .A2(new_n277), .B1(new_n762), .B2(new_n810), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n771), .A2(new_n391), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n786), .A2(G77), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n789), .B2(new_n201), .ZN(new_n1091));
  INV_X1    g0891(.A(G143), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n780), .A2(new_n208), .B1(new_n775), .B2(new_n1092), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1091), .A2(new_n1093), .A3(new_n258), .A4(new_n826), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1088), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(KEYINPUT113), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n808), .A2(G311), .B1(G317), .B2(new_n758), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT52), .Z(new_n1099));
  NAND2_X1  g0899(.A1(new_n771), .A2(G294), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n821), .A2(new_n780), .B1(new_n775), .B2(new_n801), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n374), .B(new_n1101), .C1(G107), .C2(new_n815), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n786), .A2(G116), .B1(G303), .B2(new_n788), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1096), .A2(KEYINPUT113), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1097), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1084), .B(new_n1085), .C1(new_n752), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n737), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1081), .A2(new_n1109), .ZN(G390));
  AOI21_X1  g0910(.A(new_n871), .B1(new_n714), .B2(new_n836), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n895), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n912), .B(new_n916), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n921), .A2(G330), .A3(new_n836), .A4(new_n895), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n732), .A2(new_n1116), .A3(new_n836), .A4(new_n895), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n917), .B1(new_n878), .B2(new_n895), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1113), .B(new_n1118), .C1(new_n1119), .C2(new_n913), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1113), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n845), .A2(new_n847), .B1(new_n874), .B2(new_n872), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n916), .B1(new_n1122), .B2(new_n1112), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n913), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1120), .B1(new_n1125), .B2(new_n1114), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n496), .A2(new_n612), .A3(new_n692), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n730), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n836), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1112), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1115), .A2(new_n1111), .A3(new_n1117), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1114), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n895), .B1(new_n732), .B2(new_n836), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1122), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n841), .A2(new_n715), .A3(new_n676), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n655), .B(new_n653), .C1(new_n710), .C2(new_n711), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT29), .B1(new_n1139), .B2(new_n692), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n431), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n620), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n732), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n431), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1126), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1120), .B(new_n1146), .C1(new_n1114), .C2(new_n1125), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n704), .A3(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1120), .B(new_n737), .C1(new_n1114), .C2(new_n1125), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n739), .B1(new_n275), .B2(new_n830), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G132), .A2(new_n808), .B1(new_n776), .B2(G125), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1153), .B1(new_n810), .B2(new_n785), .C1(new_n770), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n374), .B1(new_n201), .B2(new_n783), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT115), .Z(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n789), .A2(new_n962), .B1(new_n759), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n780), .A2(new_n277), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1155), .A2(new_n1157), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n770), .A2(new_n506), .B1(new_n470), .B2(new_n789), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT117), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n816), .B1(new_n465), .B2(new_n762), .C1(new_n795), .C2(new_n775), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n758), .A2(G283), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n782), .A2(new_n1090), .A3(new_n258), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1152), .B1(new_n805), .B2(new_n1170), .C1(new_n913), .C2(new_n743), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1151), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1150), .A2(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n758), .A2(G125), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n277), .B2(new_n785), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1154), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G128), .A2(new_n808), .B1(new_n781), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n817), .B2(new_n789), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G137), .C2(new_n771), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT59), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n776), .A2(G124), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n815), .C2(G159), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n770), .A2(new_n363), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G97), .A2(new_n788), .B1(new_n758), .B2(G116), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n786), .A2(G68), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n374), .A2(G41), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1055), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n783), .A2(new_n378), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n762), .A2(new_n470), .B1(new_n775), .B2(new_n792), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1187), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n329), .B1(G33), .B2(G41), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1196), .C1(new_n1190), .C2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n752), .B1(new_n1186), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n739), .B1(new_n201), .B2(new_n830), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n675), .A2(new_n290), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT118), .Z(new_n1203));
  XOR2_X1   g1003(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n302), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n614), .B1(new_n294), .B2(new_n295), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1204), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1203), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1201), .B1(new_n1212), .B2(new_n742), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT119), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n934), .B2(new_n717), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT119), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1208), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1203), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(new_n1220), .B2(new_n1209), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n923), .B1(new_n912), .B2(new_n929), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(G330), .C1(new_n1222), .C2(new_n925), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1215), .A2(KEYINPUT120), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT121), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n896), .A2(new_n918), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n1223), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n896), .A2(new_n918), .A3(KEYINPUT121), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT120), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1225), .A2(new_n1226), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1213), .B1(new_n1230), .B2(new_n737), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1149), .A2(new_n1145), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n919), .A2(new_n1223), .A3(new_n1215), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1226), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n704), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1230), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(G375));
  NOR2_X1   g1040(.A1(new_n1146), .A2(new_n1037), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1132), .A2(new_n1114), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n878), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n736), .B1(new_n1244), .B2(new_n1133), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1112), .A2(new_n742), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n771), .A2(G150), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n258), .B(new_n1192), .C1(new_n788), .C2(new_n1177), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n786), .A2(G50), .B1(G132), .B2(new_n758), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n780), .A2(new_n810), .B1(new_n775), .B2(new_n1158), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G137), .B2(new_n808), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n771), .A2(G107), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n374), .B(new_n1059), .C1(G77), .C2(new_n815), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G116), .A2(new_n788), .B1(new_n758), .B2(G294), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n762), .A2(new_n792), .B1(new_n775), .B2(new_n800), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G97), .B2(new_n781), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n805), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n739), .B(new_n1259), .C1(new_n208), .C2(new_n830), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1246), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT122), .B1(new_n1245), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1137), .A2(new_n737), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT122), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1261), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1242), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(G381));
  NOR3_X1   g1069(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1270));
  INV_X1    g1070(.A(G390), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1268), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1272), .ZN(G407));
  AOI21_X1  g1073(.A(new_n1041), .B1(new_n1126), .B2(new_n1147), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1172), .B1(new_n1274), .B2(new_n1149), .ZN(new_n1275));
  INV_X1    g1075(.A(G343), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(G213), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT123), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(G375), .C2(new_n1279), .ZN(G409));
  OAI211_X1 g1080(.A(G390), .B(new_n973), .C1(new_n1009), .C2(new_n1039), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(G396), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1271), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1281), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1288), .A3(new_n1283), .A4(new_n1281), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G378), .B(new_n1231), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1213), .B1(new_n1293), .B2(new_n737), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1232), .A2(new_n1230), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1037), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1275), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1278), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1041), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n865), .B(new_n620), .C1(new_n431), .C2(new_n1143), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(new_n1244), .A3(KEYINPUT60), .A4(new_n1133), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1302), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1302), .A2(new_n1303), .A3(new_n1305), .A4(KEYINPUT124), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1267), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1308), .A2(G384), .A3(new_n1267), .A4(new_n1309), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .A4(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1312), .A2(new_n1319), .A3(new_n1314), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1278), .A2(G2897), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1319), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1322), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1278), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1317), .B(new_n1318), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1327), .B2(new_n1316), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1291), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1332), .B1(new_n1324), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1327), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT61), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(new_n1316), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1327), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1336), .A2(new_n1290), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1331), .A2(new_n1341), .ZN(G405));
  NAND2_X1  g1142(.A1(new_n1295), .A2(new_n1233), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1041), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G378), .B1(new_n1345), .B2(new_n1231), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1292), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1289), .ZN(new_n1349));
  AOI22_X1  g1149(.A1(new_n1282), .A2(new_n1283), .B1(new_n1285), .B2(new_n1281), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1348), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1275), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1292), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1287), .A2(new_n1289), .A3(new_n1353), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1351), .A2(new_n1316), .A3(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1316), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


