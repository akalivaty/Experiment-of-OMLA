//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(G119), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT70), .A2(G128), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .A4(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(G119), .A3(new_n206), .ZN(new_n209));
  INV_X1    g023(.A(new_n202), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(KEYINPUT24), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n209), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n193), .A2(KEYINPUT74), .A3(new_n194), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n198), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n188), .A2(new_n190), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n194), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT75), .B(G110), .Z(new_n222));
  AND3_X1   g036(.A1(new_n203), .A2(new_n207), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n214), .B1(new_n209), .B2(new_n210), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n221), .B(new_n197), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT77), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT22), .B(G137), .Z(new_n232));
  OR2_X1    g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(KEYINPUT78), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n225), .A3(KEYINPUT76), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n218), .A2(new_n225), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT79), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n218), .A2(new_n225), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G217), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(G234), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G902), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n239), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n239), .A2(new_n245), .A3(KEYINPUT81), .A4(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n248), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n239), .A2(new_n245), .A3(new_n247), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT25), .ZN(new_n261));
  AOI211_X1 g075(.A(KEYINPUT82), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n259), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n261), .A3(new_n248), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G237), .A2(G953), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n269), .A2(G143), .A3(G214), .ZN(new_n270));
  AOI21_X1  g084(.A(G143), .B1(new_n269), .B2(G214), .ZN(new_n271));
  OAI21_X1  g085(.A(G131), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(G214), .ZN(new_n273));
  INV_X1    g087(.A(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n269), .A2(G143), .A3(G214), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT17), .B(G131), .C1(new_n270), .C2(new_n271), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n198), .A2(new_n217), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G113), .B(G122), .ZN(new_n285));
  INV_X1    g099(.A(G104), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT18), .A2(G131), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n275), .A2(new_n277), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n275), .B2(new_n277), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n219), .A2(KEYINPUT90), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n188), .A2(new_n190), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(G146), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n221), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT93), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n282), .A2(new_n283), .B1(new_n296), .B2(new_n291), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n287), .ZN(new_n302));
  INV_X1    g116(.A(new_n197), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n272), .B2(new_n278), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(KEYINPUT19), .A3(new_n294), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n220), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n194), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n297), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n304), .A2(new_n309), .B1(new_n291), .B2(new_n296), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n287), .B1(new_n314), .B2(KEYINPUT92), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n299), .A2(new_n302), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G475), .A2(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT94), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT20), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n313), .ZN(new_n320));
  AND4_X1   g134(.A1(new_n301), .A2(new_n284), .A3(new_n287), .A4(new_n297), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n301), .B1(new_n300), .B2(new_n287), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n324));
  INV_X1    g138(.A(new_n318), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n229), .A2(G952), .ZN(new_n328));
  INV_X1    g142(.A(G234), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(G902), .B(G953), .C1(new_n329), .C2(new_n330), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT96), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT21), .B(G898), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n321), .A2(new_n322), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n300), .A2(new_n287), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n247), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G475), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT15), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n205), .A2(G143), .A3(new_n206), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n274), .A2(G128), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G134), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n351), .B2(new_n349), .ZN(new_n354));
  XNOR2_X1  g168(.A(G116), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT95), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(G107), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(G107), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n353), .B(new_n354), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G116), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT14), .A3(G122), .ZN(new_n361));
  XOR2_X1   g175(.A(G116), .B(G122), .Z(new_n362));
  OAI211_X1 g176(.A(G107), .B(new_n361), .C1(new_n362), .C2(KEYINPUT14), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n348), .A2(new_n349), .ZN(new_n364));
  OAI221_X1 g178(.A(new_n363), .B1(G107), .B2(new_n356), .C1(new_n364), .C2(new_n350), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT83), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n367), .A2(new_n246), .A3(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n359), .B2(new_n365), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n247), .B(new_n345), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n359), .A2(new_n365), .ZN(new_n374));
  INV_X1    g188(.A(new_n368), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n369), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n345), .B1(new_n377), .B2(new_n247), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n327), .A2(new_n338), .A3(new_n342), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT97), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n319), .A2(new_n326), .B1(new_n341), .B2(G475), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n338), .A4(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G472), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT71), .A3(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n360), .A2(G119), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT2), .B(G113), .Z(new_n392));
  INV_X1    g206(.A(KEYINPUT71), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n360), .B2(G119), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT72), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n389), .A3(new_n390), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT2), .B(G113), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n194), .A2(KEYINPUT65), .A3(G143), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n274), .B2(G146), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n274), .A2(G146), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT0), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n200), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n408), .A3(new_n200), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n194), .A2(G143), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n274), .A2(G146), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n407), .A2(new_n413), .B1(new_n416), .B2(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT11), .A2(G134), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT67), .B1(new_n418), .B2(G137), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n420));
  INV_X1    g234(.A(G137), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT11), .A4(G134), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT11), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT66), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT11), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n425), .A2(new_n427), .B1(new_n349), .B2(G137), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n349), .A2(G137), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n423), .B(new_n276), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n429), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n421), .A2(G134), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n276), .B1(new_n435), .B2(new_n423), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n417), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n205), .A2(new_n206), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT1), .B1(new_n274), .B2(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n407), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT1), .ZN(new_n442));
  AND4_X1   g256(.A1(new_n442), .A2(new_n414), .A3(new_n415), .A4(G128), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n434), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n446), .A3(KEYINPUT69), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(G131), .C1(KEYINPUT69), .C2(new_n432), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n448), .A3(new_n430), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n449), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n437), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT68), .B(new_n417), .C1(new_n431), .C2(new_n436), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n402), .B(new_n450), .C1(new_n455), .C2(KEYINPUT30), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT31), .ZN(new_n457));
  INV_X1    g271(.A(new_n402), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n437), .A3(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n269), .A2(G210), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT27), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT26), .B(G101), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n456), .A2(new_n457), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n457), .B1(new_n456), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n425), .A2(new_n427), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n429), .B1(new_n472), .B2(new_n446), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n419), .A2(new_n422), .ZN(new_n474));
  OAI21_X1  g288(.A(G131), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n430), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT68), .B1(new_n476), .B2(new_n417), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n449), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n402), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n479), .B2(new_n459), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n459), .A2(new_n470), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n465), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(KEYINPUT32), .B(new_n387), .C1(new_n469), .C2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT32), .ZN(new_n485));
  INV_X1    g299(.A(new_n468), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n456), .A2(new_n457), .A3(new_n466), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n488), .B2(new_n386), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G472), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n481), .A2(new_n464), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n437), .A2(new_n449), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n402), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n459), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n464), .B1(new_n456), .B2(new_n459), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n460), .B1(new_n478), .B2(new_n402), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n481), .B(new_n464), .C1(new_n503), .C2(new_n470), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n504), .A3(new_n493), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n505), .B2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n504), .A3(new_n507), .A4(new_n493), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n491), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n268), .B(new_n385), .C1(new_n490), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G214), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G210), .B1(G237), .B2(G902), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  MUX2_X1   g328(.A(new_n417), .B(new_n445), .S(new_n189), .Z(new_n515));
  INV_X1    g329(.A(G224), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G953), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n515), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT3), .B1(new_n286), .B2(G107), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT3), .ZN(new_n523));
  INV_X1    g337(.A(G107), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(G104), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n286), .A2(G107), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT84), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(G101), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G101), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n522), .A2(new_n525), .A3(new_n532), .A4(new_n526), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n533), .A2(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n532), .A2(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n402), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G122), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n524), .A2(G104), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n286), .A2(G107), .ZN(new_n541));
  OAI21_X1  g355(.A(G101), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT5), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n388), .A3(G116), .ZN(new_n546));
  OAI211_X1 g360(.A(G113), .B(new_n546), .C1(new_n397), .C2(new_n545), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n400), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n538), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n539), .B1(new_n538), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n521), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n521), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n518), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT7), .B1(new_n516), .B2(G953), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT89), .B1(new_n445), .B2(G125), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n417), .A2(new_n189), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n445), .A2(KEYINPUT89), .A3(G125), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n539), .B(KEYINPUT8), .ZN(new_n562));
  INV_X1    g376(.A(new_n548), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n544), .B1(new_n400), .B2(new_n547), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n515), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n561), .A2(new_n549), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n247), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n514), .B1(new_n555), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  INV_X1    g385(.A(new_n551), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n549), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n553), .B1(new_n573), .B2(new_n521), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n571), .B(new_n513), .C1(new_n574), .C2(new_n518), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n512), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(G469), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  INV_X1    g393(.A(G227), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n579), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n439), .A2(G128), .B1(new_n414), .B2(new_n415), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n443), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n586), .B2(new_n543), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n415), .A2(KEYINPUT65), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n414), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(new_n403), .B1(new_n438), .B2(new_n439), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT10), .B1(new_n590), .B2(new_n443), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n591), .B2(new_n543), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n531), .A2(new_n534), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n537), .A2(new_n417), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n594), .A2(KEYINPUT85), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT85), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n537), .A2(new_n417), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n535), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n593), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n476), .ZN(new_n601));
  INV_X1    g415(.A(new_n476), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n602), .B(new_n593), .C1(new_n596), .C2(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n583), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n441), .A2(new_n543), .A3(new_n444), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n543), .B2(new_n586), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n476), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(KEYINPUT12), .A3(new_n476), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n603), .A2(new_n611), .A3(new_n583), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n578), .B(new_n247), .C1(new_n604), .C2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT86), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT85), .B1(new_n594), .B2(new_n595), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n598), .A2(new_n597), .A3(new_n535), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n476), .B(new_n592), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n617), .B2(new_n582), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n603), .A2(KEYINPUT86), .A3(new_n583), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n601), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n583), .B1(new_n603), .B2(new_n611), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n578), .B1(new_n623), .B2(new_n247), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT87), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n613), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n592), .B1(new_n615), .B2(new_n616), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n602), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n582), .B1(new_n627), .B2(new_n602), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(KEYINPUT86), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n621), .B1(new_n630), .B2(new_n618), .ZN(new_n631));
  OAI21_X1  g445(.A(G469), .B1(new_n631), .B2(G902), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n576), .B(new_n577), .C1(new_n626), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n510), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT98), .B(G101), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  INV_X1    g451(.A(new_n576), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n327), .A2(new_n342), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n377), .A2(KEYINPUT33), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n376), .A2(new_n641), .A3(new_n369), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(G478), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n377), .A2(new_n343), .A3(new_n247), .ZN(new_n644));
  NAND2_X1  g458(.A1(G478), .A2(G902), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n639), .A2(new_n647), .A3(new_n338), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT99), .B1(new_n638), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n382), .A2(new_n646), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n576), .A4(new_n338), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n577), .ZN(new_n654));
  INV_X1    g468(.A(new_n613), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n632), .B2(KEYINPUT87), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n624), .A2(new_n625), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n267), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n263), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n488), .A2(new_n247), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n488), .A2(new_n386), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n653), .A2(new_n658), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT100), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT34), .B(G104), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  NOR2_X1   g485(.A1(new_n639), .A2(new_n379), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n576), .A3(new_n338), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n658), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT35), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  INV_X1    g493(.A(KEYINPUT36), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n235), .B2(new_n236), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n228), .A2(new_n238), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n249), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n265), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n381), .B2(new_n384), .ZN(new_n689));
  INV_X1    g503(.A(new_n666), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n658), .A3(new_n690), .A4(new_n576), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  OAI21_X1  g507(.A(new_n493), .B1(new_n480), .B2(new_n492), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT73), .B1(new_n694), .B2(new_n501), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n508), .A3(new_n499), .ZN(new_n696));
  OAI22_X1  g510(.A1(new_n696), .A2(new_n491), .B1(new_n484), .B2(new_n489), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n658), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n331), .B1(new_n334), .B2(G900), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n639), .A2(new_n379), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n576), .A3(new_n687), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XNOR2_X1  g518(.A(new_n699), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n658), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT104), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n706), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n665), .A2(KEYINPUT32), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n488), .A2(new_n485), .A3(new_n386), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n456), .A2(new_n459), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n465), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n247), .B1(new_n497), .B2(new_n464), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n687), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n570), .A2(new_n575), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT38), .Z(new_n725));
  NOR4_X1   g539(.A1(new_n725), .A2(new_n512), .A3(new_n379), .A4(new_n382), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n709), .A2(new_n712), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G143), .ZN(G45));
  NOR3_X1   g542(.A1(new_n382), .A2(new_n646), .A3(new_n700), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n576), .A3(new_n687), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n698), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  NAND3_X1  g546(.A1(new_n695), .A2(new_n508), .A3(new_n499), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n713), .A2(new_n714), .B1(new_n733), .B2(G472), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n662), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n247), .B1(new_n604), .B2(new_n612), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n577), .A3(new_n613), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n737), .A2(KEYINPUT105), .A3(new_n577), .A4(new_n613), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n653), .A2(new_n735), .A3(KEYINPUT106), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n697), .A2(new_n268), .A3(new_n740), .A4(new_n741), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n649), .A2(new_n652), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NOR2_X1   g565(.A1(new_n746), .A2(new_n673), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n360), .ZN(G18));
  NAND3_X1  g567(.A1(new_n740), .A2(new_n576), .A3(new_n741), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n740), .A2(KEYINPUT107), .A3(new_n576), .A4(new_n741), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n697), .A3(new_n689), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  NAND3_X1  g573(.A1(new_n498), .A2(KEYINPUT108), .A3(new_n481), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n470), .B1(new_n496), .B2(new_n459), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n761), .B1(new_n762), .B2(new_n482), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n763), .A3(new_n465), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n486), .A3(new_n487), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n386), .ZN(new_n766));
  AOI21_X1  g580(.A(G902), .B1(new_n469), .B2(new_n483), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n660), .B(new_n766), .C1(new_n767), .C2(new_n491), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT109), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n664), .A2(new_n770), .A3(new_n660), .A4(new_n766), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n742), .A2(new_n337), .ZN(new_n773));
  INV_X1    g587(.A(new_n379), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n639), .A2(KEYINPUT110), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n382), .B2(new_n379), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n777), .A3(new_n576), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT111), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G122), .ZN(G24));
  NAND4_X1  g598(.A1(new_n664), .A2(new_n729), .A3(new_n687), .A4(new_n766), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n756), .A2(new_n757), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  NAND2_X1  g602(.A1(new_n265), .A2(new_n266), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n734), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(G902), .B1(new_n620), .B2(new_n622), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n613), .B1(new_n791), .B2(new_n578), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n570), .A2(new_n575), .A3(new_n511), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n793), .A3(new_n577), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n790), .A2(KEYINPUT42), .A3(new_n729), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n697), .A2(new_n794), .A3(new_n268), .A4(new_n729), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  NAND3_X1  g616(.A1(new_n735), .A2(new_n701), .A3(new_n794), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G134), .ZN(G36));
  OR3_X1    g618(.A1(new_n639), .A2(KEYINPUT43), .A3(new_n646), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n647), .A2(new_n382), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT43), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n690), .A2(new_n688), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT44), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(new_n811), .A3(KEYINPUT44), .A4(new_n810), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n793), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n578), .B1(new_n623), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n817), .B2(new_n623), .ZN(new_n819));
  NAND2_X1  g633(.A1(G469), .A2(G902), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT46), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT114), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n613), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n819), .A2(KEYINPUT46), .A3(new_n820), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT113), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n577), .B(new_n705), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  AND2_X1   g646(.A1(new_n729), .A2(new_n793), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n734), .A2(new_n833), .A3(new_n662), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n577), .B1(new_n827), .B2(new_n829), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT47), .B(new_n577), .C1(new_n827), .C2(new_n829), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(new_n187), .ZN(G42));
  OAI211_X1 g654(.A(new_n658), .B(new_n697), .C1(new_n702), .C2(new_n730), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n576), .A2(new_n775), .A3(new_n777), .A4(new_n699), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n654), .B1(new_n632), .B2(new_n613), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n721), .A3(new_n688), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n787), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n787), .A2(new_n841), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n746), .A2(new_n673), .B1(new_n510), .B2(new_n634), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n783), .A2(new_n853), .A3(new_n749), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n664), .A2(new_n687), .A3(new_n766), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n794), .A4(new_n729), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n843), .A2(new_n793), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n785), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n793), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n382), .A2(new_n379), .A3(new_n699), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n861), .A2(new_n688), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n658), .A3(new_n697), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n803), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n796), .A2(new_n798), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n865), .B1(new_n869), .B2(new_n795), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n638), .A2(new_n648), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n667), .A2(new_n658), .A3(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n675), .A2(new_n758), .A3(new_n691), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n851), .A2(new_n854), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n852), .B1(new_n748), .B2(new_n744), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n873), .A3(new_n783), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n860), .A2(new_n803), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n801), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n787), .A2(new_n841), .A3(new_n846), .A4(new_n844), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n874), .B(new_n875), .C1(new_n883), .C2(KEYINPUT53), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT117), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT117), .B1(new_n877), .B2(new_n879), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n848), .A3(new_n850), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n884), .B1(new_n890), .B2(new_n875), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n662), .A2(new_n331), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n742), .A2(new_n861), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n722), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n639), .A3(new_n647), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n808), .A2(new_n331), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n893), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n855), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n896), .A2(new_n772), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n743), .A2(new_n512), .A3(new_n725), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n899), .A2(KEYINPUT50), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT50), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n737), .A2(new_n613), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n654), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n837), .A2(new_n838), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n899), .A2(new_n793), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT119), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT51), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n897), .A2(new_n790), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT48), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n756), .A3(new_n757), .ZN(new_n913));
  INV_X1    g727(.A(new_n650), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n913), .B(new_n328), .C1(new_n914), .C2(new_n894), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n908), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n901), .A2(new_n902), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n898), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n909), .A2(KEYINPUT120), .A3(KEYINPUT51), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n910), .B(new_n916), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n891), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n904), .B(KEYINPUT49), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n806), .A2(new_n789), .A3(new_n512), .A4(new_n654), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n722), .A2(new_n926), .A3(new_n725), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n229), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n874), .B1(new_n883), .B2(KEYINPUT53), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(G902), .ZN(new_n934));
  INV_X1    g748(.A(G210), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n574), .B(new_n518), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT121), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n936), .A2(new_n942), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n941), .B2(new_n943), .ZN(G51));
  NOR2_X1   g758(.A1(new_n934), .A2(new_n819), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n604), .A2(new_n612), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n933), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n884), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n820), .B(KEYINPUT57), .Z(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n947), .B2(new_n884), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT122), .B1(new_n954), .B2(new_n946), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n930), .B1(new_n952), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(new_n933), .A2(G902), .ZN(new_n957));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT123), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n323), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n957), .A2(new_n959), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n930), .B1(new_n964), .B2(new_n316), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(G60));
  AND2_X1   g780(.A1(new_n640), .A2(new_n642), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n645), .B(KEYINPUT59), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n948), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n931), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n891), .A2(new_n969), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n967), .ZN(G63));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT60), .Z(new_n976));
  AND2_X1   g790(.A1(new_n933), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(new_n685), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n930), .B1(new_n977), .B2(new_n685), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n933), .A2(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n239), .A2(new_n245), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n983), .B(new_n980), .C1(new_n978), .C2(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G66));
  OAI21_X1  g801(.A(G953), .B1(new_n336), .B2(new_n516), .ZN(new_n988));
  INV_X1    g802(.A(new_n877), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(G953), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n574), .B1(G898), .B2(new_n229), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G69));
  OAI21_X1  g806(.A(new_n450), .B1(new_n455), .B2(KEYINPUT30), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n305), .A2(new_n308), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(new_n995));
  INV_X1    g809(.A(new_n839), .ZN(new_n996));
  INV_X1    g810(.A(new_n830), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n778), .A3(new_n790), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n787), .A2(new_n841), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n801), .A2(new_n803), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n996), .A2(new_n831), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n229), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n580), .A2(G900), .A3(G953), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n727), .A2(new_n1006), .A3(new_n999), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n727), .A2(new_n1009), .A3(new_n1006), .A4(new_n999), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1006), .B1(new_n727), .B2(new_n999), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n735), .B(new_n793), .C1(new_n650), .C2(new_n672), .ZN(new_n1013));
  OAI22_X1  g827(.A1(new_n816), .A2(new_n830), .B1(new_n711), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1012), .A2(new_n839), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1005), .B1(new_n1016), .B2(G953), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1004), .B1(new_n1017), .B2(new_n995), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1001), .B2(new_n877), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n716), .A2(new_n464), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n930), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n718), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1022), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1024), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n890), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n1016), .B2(new_n877), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n718), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT127), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1028), .A2(new_n1031), .A3(new_n718), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1027), .B1(new_n1030), .B2(new_n1032), .ZN(G57));
endmodule


