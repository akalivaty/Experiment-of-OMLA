//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT68), .B(G77), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AND2_X1   g0008(.A1(new_n208), .A2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G58), .A2(G232), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT67), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(KEYINPUT66), .A2(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(KEYINPUT66), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n218), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n226), .B(new_n230), .C1(KEYINPUT1), .C2(new_n215), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n242), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n219), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT70), .B1(new_n251), .B2(new_n219), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n223), .A2(new_n207), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n260), .B(KEYINPUT72), .Z(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT15), .B(G87), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G33), .A3(new_n223), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT73), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n256), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n252), .B(new_n253), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT69), .A2(G1), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT69), .A2(G1), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT69), .A2(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT69), .A2(G1), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(G13), .A3(G20), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n273), .A2(G77), .B1(new_n207), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G107), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G238), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n283), .B1(new_n284), .B2(new_n281), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n220), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n220), .A2(new_n291), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n274), .A2(new_n275), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n299), .B2(G244), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G190), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n280), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n279), .B(new_n307), .C1(G169), .C2(new_n303), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n258), .A2(G150), .ZN(new_n311));
  INV_X1    g0111(.A(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n223), .A2(G33), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n312), .B2(new_n201), .C1(new_n313), .C2(new_n257), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n256), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n277), .A2(new_n243), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n316), .C1(new_n243), .C2(new_n272), .ZN(new_n317));
  OR2_X1    g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(G1698), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G222), .ZN(new_n321));
  INV_X1    g0121(.A(G223), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n321), .B1(new_n207), .B2(new_n281), .C1(new_n285), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n288), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n295), .B1(new_n299), .B2(G226), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n317), .B1(new_n327), .B2(G169), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n306), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n317), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n317), .A2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n335), .B2(new_n341), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n310), .B(new_n332), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(new_n282), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n281), .A2(new_n350), .A3(G226), .A4(new_n282), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G232), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT76), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(G33), .A3(G97), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n296), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n292), .A2(new_n294), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n298), .B2(new_n286), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT13), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n351), .B2(new_n349), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(new_n296), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(G169), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT77), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n369), .A2(KEYINPUT77), .A3(new_n370), .A4(G169), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n368), .A3(G179), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n276), .A2(G68), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n245), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n313), .B2(new_n202), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT11), .B1(new_n382), .B2(new_n256), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n245), .B2(new_n272), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n339), .B2(new_n369), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n364), .B2(new_n368), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G232), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n362), .B1(new_n298), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n322), .A2(new_n282), .ZN(new_n398));
  INV_X1    g0198(.A(G226), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(new_n400), .C1(new_n346), .C2(new_n347), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT80), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n296), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n401), .A2(KEYINPUT80), .A3(new_n402), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  INV_X1    g0208(.A(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  INV_X1    g0210(.A(new_n257), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n277), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n272), .B2(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n318), .A2(new_n312), .A3(new_n319), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  AND2_X1   g0216(.A1(KEYINPUT78), .A2(KEYINPUT7), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT78), .A2(KEYINPUT7), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n346), .A2(new_n347), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n223), .A2(new_n421), .A3(KEYINPUT7), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n416), .B1(new_n415), .B2(new_n419), .ZN(new_n424));
  OAI21_X1  g0224(.A(G68), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G58), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n245), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G58), .A2(G68), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n258), .A2(G159), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT7), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT66), .A2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT66), .A2(G20), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n318), .A3(new_n436), .A4(new_n319), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n346), .A2(new_n347), .A3(G20), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n434), .A2(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT16), .B(new_n432), .C1(new_n440), .C2(new_n245), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n256), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n414), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n410), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n410), .B2(new_n443), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT81), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n425), .A2(new_n432), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT16), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(new_n434), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n438), .A2(new_n439), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n431), .B1(new_n453), .B2(G68), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n267), .B1(new_n454), .B2(KEYINPUT16), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n413), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n405), .A2(new_n406), .ZN(new_n457));
  INV_X1    g0257(.A(new_n397), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n457), .A2(G179), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n409), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT18), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n410), .A2(new_n443), .A3(new_n444), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n457), .A2(G190), .A3(new_n458), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n391), .B1(new_n457), .B2(new_n458), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n450), .A2(new_n455), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT17), .A4(new_n414), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n457), .A2(G190), .A3(new_n458), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n391), .B2(new_n407), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n443), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n447), .A2(new_n465), .A3(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n345), .A2(new_n395), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n277), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n270), .A2(G33), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n276), .C1(new_n254), .C2(new_n255), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(new_n478), .ZN(new_n482));
  INV_X1    g0282(.A(G33), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n435), .A2(new_n484), .A3(new_n436), .A4(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n251), .A2(new_n219), .B1(G20), .B2(new_n478), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n486), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT20), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(new_n282), .C1(new_n346), .C2(new_n347), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n492), .B(new_n493), .C1(new_n494), .C2(new_n281), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n495), .A2(new_n288), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n274), .A2(G45), .A3(new_n275), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G270), .B(new_n296), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n268), .A2(new_n269), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n498), .A2(new_n499), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n292), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(KEYINPUT86), .B(new_n491), .C1(new_n510), .C2(new_n391), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(G190), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n495), .A2(new_n288), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n508), .B1(new_n501), .B2(new_n505), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT86), .B1(new_n518), .B2(new_n491), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  OAI21_X1  g0321(.A(G179), .B1(new_n482), .B2(new_n490), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n479), .B1(new_n488), .B2(new_n489), .C1(new_n481), .C2(new_n478), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n510), .A2(KEYINPUT85), .A3(G179), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(new_n524), .A3(G169), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n517), .A2(new_n524), .A3(KEYINPUT21), .A4(G169), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n288), .B1(new_n503), .B2(new_n504), .ZN(new_n533));
  OAI211_X1 g0333(.A(G257), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(new_n282), .C1(new_n346), .C2(new_n347), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G294), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(G264), .A2(new_n533), .B1(new_n537), .B2(new_n288), .ZN(new_n538));
  AOI21_X1  g0338(.A(G169), .B1(new_n538), .B2(new_n505), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n288), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n296), .C1(new_n497), .C2(new_n500), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n505), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(G179), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n435), .B(new_n436), .C1(new_n346), .C2(new_n347), .ZN(new_n545));
  INV_X1    g0345(.A(G87), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT22), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n223), .A2(new_n281), .A3(new_n548), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n223), .A2(KEYINPUT23), .A3(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(KEYINPUT23), .A2(G107), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n554));
  OAI221_X1 g0354(.A(new_n552), .B1(KEYINPUT87), .B2(new_n553), .C1(new_n554), .C2(G20), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(KEYINPUT87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n550), .A2(new_n556), .A3(KEYINPUT87), .A4(new_n553), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n267), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n276), .A2(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n284), .B2(new_n481), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n544), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n281), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n281), .A2(G238), .A3(new_n282), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n288), .ZN(new_n573));
  INV_X1    g0373(.A(G250), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n288), .B1(new_n497), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n503), .A2(new_n290), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n306), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n435), .A2(G33), .A3(G97), .A4(new_n436), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n223), .A2(new_n281), .A3(G68), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT19), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n223), .B1(new_n546), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n256), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n277), .A2(new_n262), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n267), .A2(new_n276), .A3(new_n263), .A4(new_n480), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n572), .A2(new_n288), .B1(new_n576), .B2(new_n575), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n578), .B(new_n590), .C1(G169), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n573), .A2(new_n577), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G200), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(G190), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n267), .A2(G87), .A3(new_n276), .A4(new_n480), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n587), .A2(new_n588), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n565), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(G107), .B1(new_n423), .B2(new_n424), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n284), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  XOR2_X1   g0401(.A(G97), .B(G107), .Z(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(KEYINPUT6), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n224), .B1(G77), .B2(new_n258), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n256), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n296), .C1(new_n497), .C2(new_n500), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n505), .ZN(new_n608));
  OAI211_X1 g0408(.A(G244), .B(new_n282), .C1(new_n346), .C2(new_n347), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n485), .A4(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n608), .B1(new_n288), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n485), .B(new_n613), .C1(new_n609), .C2(new_n610), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT4), .B1(new_n320), .B2(G244), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n288), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n607), .A2(new_n505), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  INV_X1    g0422(.A(G97), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n277), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n481), .B2(new_n623), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n606), .A2(new_n616), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n409), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n619), .A2(new_n620), .A3(new_n306), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n267), .B1(new_n600), .B2(new_n604), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n625), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT82), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n599), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT82), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n559), .A2(new_n560), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n564), .B1(new_n635), .B2(new_n256), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n542), .A2(new_n391), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT88), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n542), .A2(new_n639), .A3(new_n391), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n538), .A2(new_n339), .A3(new_n505), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n477), .A2(new_n532), .A3(new_n633), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n332), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n389), .B1(new_n393), .B2(new_n308), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n475), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n462), .A2(new_n464), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n343), .A2(new_n344), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n477), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n572), .A2(KEYINPUT89), .A3(new_n288), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT89), .B1(new_n572), .B2(new_n288), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n577), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n409), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n578), .A2(new_n590), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI221_X4 g0460(.A(new_n339), .B1(new_n576), .B2(new_n575), .C1(new_n572), .C2(new_n288), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n587), .A2(new_n588), .A3(new_n596), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT89), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n573), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n572), .A2(KEYINPUT89), .A3(new_n288), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n576), .B2(new_n575), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n667), .B2(new_n391), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n630), .A2(new_n625), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n629), .B1(new_n615), .B2(G169), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n660), .A2(new_n668), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n606), .A2(new_n626), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n619), .A2(new_n306), .A3(new_n620), .ZN(new_n675));
  AOI21_X1  g0475(.A(G169), .B1(new_n619), .B2(new_n620), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n598), .A2(new_n674), .A3(new_n592), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n673), .A2(new_n679), .A3(KEYINPUT90), .A4(new_n660), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n565), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n627), .A2(new_n631), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n657), .A2(G200), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n659), .A2(new_n658), .B1(new_n683), .B2(new_n663), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n643), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n678), .A2(KEYINPUT26), .B1(new_n659), .B2(new_n658), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT90), .B1(new_n687), .B2(new_n673), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n653), .B1(new_n654), .B2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n223), .A2(G13), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n270), .ZN(new_n694));
  INV_X1    g0494(.A(G213), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n692), .A2(KEYINPUT27), .A3(new_n297), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n524), .ZN(new_n700));
  MUX2_X1   g0500(.A(new_n531), .B(new_n532), .S(new_n700), .Z(new_n701));
  NOR2_X1   g0501(.A1(new_n636), .A2(new_n698), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n636), .B2(new_n642), .ZN(new_n703));
  INV_X1    g0503(.A(new_n565), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n565), .A2(new_n699), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n701), .A2(new_n707), .A3(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n531), .A2(new_n698), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n705), .A2(new_n709), .B1(new_n565), .B2(new_n699), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n698), .C1(new_n686), .C2(new_n688), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n678), .A2(new_n669), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT94), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n684), .A2(KEYINPUT26), .A3(new_n672), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n678), .A2(new_n719), .A3(new_n669), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n643), .A2(new_n660), .A3(new_n668), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n682), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n627), .A2(new_n631), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT95), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n722), .A2(new_n681), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n660), .B(KEYINPUT93), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n721), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n713), .B1(new_n729), .B2(new_n698), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n715), .A2(new_n730), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n532), .A2(new_n633), .A3(new_n644), .A4(new_n698), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n306), .B1(new_n495), .B2(new_n288), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n538), .B(new_n733), .C1(new_n515), .C2(new_n516), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n615), .A4(new_n591), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n538), .B2(new_n505), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n657), .A2(new_n517), .A3(new_n621), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n615), .A2(new_n591), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n734), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n736), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT92), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n742), .A2(KEYINPUT92), .A3(KEYINPUT31), .A4(new_n699), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n699), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n732), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n731), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G1), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n227), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G41), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n585), .A2(new_n546), .A3(new_n478), .ZN(new_n758));
  OR3_X1    g0558(.A1(new_n757), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n217), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n762));
  XNOR2_X1  g0562(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n763), .ZN(G364));
  AOI21_X1  g0564(.A(new_n754), .B1(new_n693), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n757), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n701), .B2(G330), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n701), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT96), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n249), .A2(new_n502), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n756), .A2(new_n281), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n772), .B(new_n774), .C1(new_n502), .C2(new_n218), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n756), .A2(new_n421), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n478), .B2(new_n756), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT97), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n219), .B1(G20), .B2(new_n409), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n767), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n784), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n701), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n224), .A2(new_n339), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n391), .A2(G179), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n224), .A2(new_n339), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n284), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n223), .B1(G190), .B2(new_n791), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n623), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(G20), .A3(G190), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n546), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n798), .A2(new_n800), .A3(new_n421), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n223), .A2(new_n306), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n339), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G200), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n804), .B1(new_n208), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n806), .A2(G190), .A3(new_n391), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G50), .A2(new_n811), .B1(new_n812), .B2(G58), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n339), .A3(G200), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n809), .B(new_n813), .C1(new_n245), .C2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  INV_X1    g0616(.A(new_n797), .ZN(new_n817));
  INV_X1    g0617(.A(new_n792), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n817), .B1(new_n818), .B2(G329), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT100), .Z(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G322), .B2(new_n812), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n421), .B1(new_n494), .B2(new_n801), .C1(new_n799), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n811), .B2(G326), .ZN(new_n824));
  INV_X1    g0624(.A(new_n814), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G311), .A2(new_n808), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n821), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n816), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n788), .B(new_n790), .C1(new_n785), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n771), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT101), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(G396));
  AOI22_X1  g0636(.A1(new_n808), .A2(G159), .B1(new_n812), .B2(G143), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n810), .C1(new_n839), .C2(new_n814), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  NOR2_X1   g0641(.A1(new_n797), .A2(new_n245), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n281), .B1(new_n801), .B2(new_n243), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n792), .A2(new_n844), .B1(new_n799), .B2(new_n426), .ZN(new_n845));
  NOR4_X1   g0645(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n808), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n847), .A2(new_n478), .B1(new_n494), .B2(new_n810), .ZN(new_n848));
  INV_X1    g0648(.A(new_n812), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n822), .B1(new_n850), .B2(new_n814), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G87), .A2(new_n817), .B1(new_n818), .B2(G311), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n853));
  INV_X1    g0653(.A(new_n801), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n281), .B(new_n800), .C1(G107), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n848), .A2(new_n851), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n785), .B1(new_n846), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n767), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n785), .A2(new_n782), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n202), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n280), .A2(new_n302), .A3(new_n304), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n280), .A2(new_n698), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n308), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n308), .A2(new_n699), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n859), .B(new_n862), .C1(new_n783), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n752), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n673), .A2(new_n679), .A3(new_n660), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT90), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n685), .A3(new_n680), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n868), .B1(new_n874), .B2(new_n698), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT103), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n309), .A2(new_n699), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n686), .B2(new_n688), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n870), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT104), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n870), .A3(new_n878), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n860), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n879), .A2(KEYINPUT104), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n869), .B1(new_n882), .B2(new_n883), .ZN(G384));
  XOR2_X1   g0684(.A(new_n603), .B(KEYINPUT105), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n886), .A2(G116), .A3(new_n220), .A4(new_n224), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT36), .ZN(new_n890));
  OR3_X1    g0690(.A1(new_n207), .A2(new_n217), .A3(new_n427), .ZN(new_n891));
  AOI211_X1 g0691(.A(G13), .B(new_n270), .C1(new_n891), .C2(new_n244), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n865), .A2(new_n867), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n388), .A2(new_n699), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n389), .A2(new_n394), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n388), .B(new_n699), .C1(new_n378), .C2(new_n393), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n532), .A2(new_n633), .A3(new_n644), .A4(new_n698), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT31), .B1(new_n742), .B2(new_n699), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n454), .A2(KEYINPUT16), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n414), .B1(new_n906), .B2(new_n442), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n410), .B2(new_n697), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n456), .A2(new_n468), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n410), .A2(new_n443), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n443), .A2(new_n697), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n909), .A2(new_n912), .A3(new_n913), .A4(new_n905), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n697), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI221_X4 g0716(.A(new_n904), .B1(new_n911), .B2(new_n914), .C1(new_n476), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n914), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n470), .A2(new_n474), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n443), .B(new_n697), .C1(new_n649), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n898), .B(new_n903), .C1(new_n917), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n649), .B2(KEYINPUT81), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n915), .B1(new_n925), .B2(new_n465), .ZN(new_n926));
  INV_X1    g0726(.A(new_n918), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n910), .B1(new_n927), .B2(new_n905), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n904), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n476), .A2(new_n916), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n911), .A2(new_n914), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n896), .A2(new_n897), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n934), .A2(new_n903), .A3(new_n868), .ZN(new_n935));
  AOI22_X1  g0735(.A1(KEYINPUT40), .A2(new_n924), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n477), .A2(new_n903), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(G330), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n917), .B2(new_n923), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n378), .A2(new_n388), .A3(new_n698), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n650), .A2(new_n697), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n878), .A2(new_n867), .B1(new_n896), .B2(new_n897), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n929), .A2(new_n932), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n477), .B1(new_n715), .B2(new_n730), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n653), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n942), .A2(new_n956), .B1(new_n270), .B2(new_n693), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n942), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n893), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI21_X1  g0759(.A(new_n684), .B1(new_n597), .B2(new_n698), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n658), .A2(new_n659), .A3(new_n662), .A4(new_n699), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n724), .B(new_n726), .C1(new_n670), .C2(new_n698), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n672), .A2(new_n699), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT106), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT106), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT42), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n631), .B1(new_n968), .B2(new_n565), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n698), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT107), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n965), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n963), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(KEYINPUT108), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n708), .A2(new_n971), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n981), .A2(new_n964), .A3(new_n963), .A4(new_n983), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n991), .B(new_n965), .C1(new_n981), .C2(new_n983), .ZN(new_n992));
  INV_X1    g0792(.A(new_n989), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n711), .B2(new_n970), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n971), .A2(new_n710), .A3(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n971), .B2(new_n710), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n998), .A2(new_n1002), .A3(new_n708), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n708), .B1(new_n998), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n709), .B1(new_n705), .B2(new_n706), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n967), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n701), .A2(G330), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT109), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1007), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n753), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n757), .B(KEYINPUT41), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n765), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n990), .A2(new_n994), .A3(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n786), .B1(new_n227), .B2(new_n262), .C1(new_n774), .C2(new_n238), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(new_n767), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT110), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n817), .A2(G97), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n818), .A2(G317), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n421), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n811), .A2(G311), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT46), .B1(new_n801), .B2(new_n478), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n801), .A2(KEYINPUT46), .A3(new_n478), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n799), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1023), .A2(new_n1024), .B1(new_n1025), .B2(G107), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1026), .C1(new_n822), .C2(new_n814), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n812), .A2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n1018), .B2(new_n1021), .C1(new_n847), .C2(new_n850), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G143), .A2(new_n811), .B1(new_n812), .B2(G150), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n793), .B2(new_n814), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n281), .B1(new_n801), .B2(new_n426), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n799), .A2(new_n245), .B1(new_n797), .B2(new_n207), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G137), .C2(new_n818), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n847), .B2(new_n243), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1027), .A2(new_n1029), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT47), .Z(new_n1037));
  INV_X1    g0837(.A(new_n785), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1017), .B1(new_n789), .B2(new_n962), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1015), .A2(new_n1039), .ZN(G387));
  NOR2_X1   g0840(.A1(new_n235), .A2(new_n502), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n411), .A2(KEYINPUT50), .A3(new_n243), .ZN(new_n1042));
  AOI21_X1  g0842(.A(KEYINPUT50), .B1(new_n411), .B2(new_n243), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n758), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n774), .B(new_n1041), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n776), .A2(new_n758), .B1(new_n284), .B2(new_n756), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1046), .B1(KEYINPUT112), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT112), .B2(new_n1048), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n860), .B1(new_n1050), .B2(new_n786), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n707), .B2(new_n789), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n808), .B1(new_n825), .B2(new_n411), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n799), .A2(new_n262), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G150), .B2(new_n818), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n421), .B1(new_n854), .B2(new_n208), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n1019), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n812), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1053), .B(new_n1058), .C1(new_n793), .C2(new_n810), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n281), .B1(new_n818), .B2(G326), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n799), .A2(new_n850), .B1(new_n822), .B2(new_n801), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G311), .A2(new_n825), .B1(new_n811), .B2(G322), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n808), .A2(G303), .B1(new_n812), .B2(G317), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1060), .B1(new_n478), .B2(new_n797), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1059), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1038), .B1(new_n1071), .B2(KEYINPUT113), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1052), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1011), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT111), .B1(new_n1075), .B2(new_n765), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT111), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1011), .A2(new_n1077), .A3(new_n766), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n753), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1011), .A2(new_n731), .A3(new_n752), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n757), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1079), .A2(new_n1082), .ZN(G393));
  INV_X1    g0883(.A(new_n1005), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n757), .B1(new_n1084), .B2(new_n1081), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1081), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1005), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n970), .A2(new_n789), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n773), .A2(new_n242), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n787), .B1(new_n756), .B2(G97), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n860), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G150), .A2(new_n811), .B1(new_n812), .B2(G159), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT115), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT51), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n799), .A2(new_n202), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n281), .B1(new_n245), .B2(new_n801), .C1(new_n797), .C2(new_n546), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(G143), .C2(new_n818), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n243), .B2(new_n814), .C1(new_n847), .C2(new_n257), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1095), .B2(KEYINPUT51), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G317), .A2(new_n811), .B1(new_n812), .B2(G311), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  AOI22_X1  g0903(.A1(new_n818), .A2(G322), .B1(G283), .B2(new_n854), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G294), .A2(new_n808), .B1(new_n825), .B2(G303), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n281), .B(new_n798), .C1(G116), .C2(new_n1025), .ZN(new_n1108));
  AND4_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1096), .A2(new_n1101), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1090), .B(new_n1093), .C1(new_n1038), .C2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1084), .B2(new_n765), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1088), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n944), .A2(new_n945), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n782), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n861), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n767), .B1(new_n411), .B2(new_n1117), .ZN(new_n1118));
  OR3_X1    g0918(.A1(new_n1097), .A2(new_n281), .A3(new_n802), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n842), .B1(G294), .B2(new_n818), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT118), .Z(new_n1121));
  AOI22_X1  g0921(.A1(G107), .A2(new_n825), .B1(new_n812), .B2(G116), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n850), .C2(new_n810), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1119), .B(new_n1123), .C1(G97), .C2(new_n808), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(KEYINPUT119), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(KEYINPUT119), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n847), .A2(new_n1127), .B1(new_n838), .B2(new_n814), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G132), .B2(new_n812), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n811), .A2(G128), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT53), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n854), .B2(G150), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1132), .A2(new_n421), .A3(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n797), .A2(new_n243), .B1(new_n799), .B2(new_n793), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G125), .B2(new_n818), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1129), .A2(new_n1130), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1125), .A2(new_n1126), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1138), .B2(new_n785), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT117), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n950), .B2(new_n947), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n866), .B1(new_n874), .B2(new_n877), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n934), .ZN(new_n1144));
  OAI211_X1 g0944(.A(KEYINPUT117), .B(new_n946), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1115), .A3(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n868), .B(G330), .C1(new_n732), .C2(new_n750), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n1144), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n729), .A2(new_n698), .A3(new_n865), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n867), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n934), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n946), .B1(new_n917), .B2(new_n923), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1148), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n766), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n941), .B1(new_n899), .B2(new_n902), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n898), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1144), .B1(new_n1149), .B2(new_n867), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1152), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1146), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1140), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n477), .A2(new_n1157), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n954), .A2(new_n653), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1147), .A2(new_n1144), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1143), .B1(new_n1169), .B2(new_n1158), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n934), .B1(new_n1157), .B2(new_n868), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1148), .A2(new_n1150), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1168), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1147), .A2(new_n1144), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1159), .B2(new_n1152), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n946), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1176), .A2(new_n1141), .B1(new_n944), .B2(new_n945), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n1145), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1173), .B1(new_n1162), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1170), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1150), .A2(new_n1171), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1174), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1167), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1160), .B1(new_n1177), .B2(new_n1145), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1155), .C1(new_n1184), .C2(new_n1158), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1179), .A2(new_n1185), .A3(new_n757), .ZN(new_n1186));
  OAI211_X1 g0986(.A(KEYINPUT120), .B(new_n1140), .C1(new_n1156), .C2(new_n1162), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1165), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT121), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT121), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1165), .A2(new_n1186), .A3(new_n1190), .A4(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(G378));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n652), .A2(new_n332), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n317), .A2(new_n697), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT40), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n951), .A2(new_n935), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n928), .B1(new_n476), .B2(new_n916), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n923), .B1(new_n1201), .B2(KEYINPUT38), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n934), .A2(new_n903), .A3(new_n868), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT40), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n941), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1205), .A2(new_n953), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n953), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1198), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n948), .B(new_n952), .C1(new_n936), .C2(new_n941), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1196), .B(new_n1197), .Z(new_n1210));
  NAND2_X1  g1010(.A1(new_n1205), .A2(new_n953), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1193), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1185), .A2(new_n1168), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n760), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1210), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1162), .A2(new_n1178), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1172), .A2(new_n1170), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1167), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1193), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1215), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1210), .A2(new_n782), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n767), .B1(G50), .B2(new_n1117), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G33), .A2(G41), .ZN(new_n1228));
  INV_X1    g1028(.A(G41), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G50), .B(new_n1228), .C1(new_n421), .C2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n797), .A2(new_n426), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G283), .B2(new_n818), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G41), .B(new_n281), .C1(new_n854), .C2(new_n208), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n245), .C2(new_n799), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G107), .B2(new_n812), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n263), .A2(new_n808), .B1(new_n811), .B2(G116), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n623), .C2(new_n814), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1230), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n799), .A2(new_n839), .B1(new_n801), .B2(new_n1127), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G125), .A2(new_n811), .B1(new_n812), .B2(G128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n838), .B2(new_n847), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G132), .C2(new_n825), .ZN(new_n1243));
  XOR2_X1   g1043(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1228), .B1(new_n797), .B2(new_n793), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G124), .B2(new_n818), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1239), .B1(new_n1238), .B2(new_n1237), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1227), .B1(new_n1250), .B2(new_n785), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1225), .A2(new_n766), .B1(new_n1226), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1224), .A2(new_n1252), .ZN(G375));
  NAND2_X1  g1053(.A1(new_n1220), .A2(new_n1167), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1013), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1173), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1144), .A2(new_n782), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n767), .B1(G68), .B2(new_n1117), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n281), .B(new_n1054), .C1(G97), .C2(new_n854), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n202), .B2(new_n797), .C1(new_n494), .C2(new_n792), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G107), .B2(new_n808), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G116), .A2(new_n825), .B1(new_n812), .B2(G283), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n822), .C2(new_n810), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n844), .A2(new_n810), .B1(new_n814), .B2(new_n1127), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G137), .B2(new_n812), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT123), .Z(new_n1266));
  AOI211_X1 g1066(.A(new_n421), .B(new_n1231), .C1(G159), .C2(new_n854), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n818), .A2(G128), .B1(new_n1025), .B2(G50), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(new_n847), .C2(new_n839), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1263), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1258), .B1(new_n1270), .B2(new_n785), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1221), .A2(new_n766), .B1(new_n1257), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1256), .A2(new_n1272), .ZN(G381));
  AND3_X1   g1073(.A1(new_n1113), .A2(new_n1015), .A3(new_n1039), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n766), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1163), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1186), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1283), .A2(G384), .A3(G381), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1274), .A2(new_n1278), .A3(new_n1281), .A4(new_n1284), .ZN(G407));
  NOR2_X1   g1085(.A1(new_n695), .A2(G343), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1278), .A2(new_n1281), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G407), .A2(G213), .A3(new_n1287), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G393), .A2(G396), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1282), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1113), .B1(new_n1039), .B2(new_n1015), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1292), .C1(new_n1274), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1113), .A2(new_n1015), .A3(new_n1039), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1283), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT125), .B1(new_n1291), .B2(new_n1282), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n882), .A2(new_n883), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1220), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n757), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1173), .A2(KEYINPUT60), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1254), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1272), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1301), .B(new_n869), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1304), .A2(new_n1254), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1272), .C1(new_n1308), .C2(new_n1303), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1286), .A2(G2897), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(G2897), .A3(new_n1286), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1225), .A2(new_n1214), .A3(new_n1255), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1280), .B1(new_n1252), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(G378), .B2(new_n1278), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1313), .B(new_n1314), .C1(new_n1317), .C2(new_n1286), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1317), .A2(new_n1286), .A3(new_n1310), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1318), .B(new_n1319), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G378), .A2(new_n1278), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1286), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1311), .A3(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1327), .A2(KEYINPUT62), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1300), .B1(new_n1322), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT63), .B1(new_n1320), .B2(KEYINPUT124), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1300), .A2(KEYINPUT61), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1330), .A2(new_n1333), .A3(new_n1334), .A4(new_n1318), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1281), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1323), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1311), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1338), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1337), .A2(new_n1339), .A3(new_n1323), .A4(new_n1311), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1300), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1344), .B(new_n1345), .ZN(G402));
endmodule


