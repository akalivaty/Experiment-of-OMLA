//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT68), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n209), .B2(new_n204), .ZN(new_n210));
  XOR2_X1   g009(.A(G127gat), .B(G134gat), .Z(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(new_n204), .B2(new_n207), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT23), .B1(new_n218), .B2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n221), .C1(G169gat), .C2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  AND4_X1   g022(.A1(KEYINPUT25), .A2(new_n219), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT65), .A3(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n228), .A2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n227), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n226), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n241), .A2(new_n228), .A3(new_n229), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  NOR3_X1   g043(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n218), .B1(new_n246), .B2(new_n223), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT27), .B(G183gat), .ZN(new_n248));
  INV_X1    g047(.A(G190gat), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(KEYINPUT28), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT28), .B1(new_n248), .B2(new_n249), .ZN(new_n251));
  OAI221_X1 g050(.A(new_n225), .B1(new_n245), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n238), .B1(new_n237), .B2(new_n243), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n217), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n253), .A2(new_n217), .A3(new_n254), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n217), .C1(new_n253), .C2(new_n254), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n202), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT32), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g062(.A(new_n259), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n237), .A2(new_n243), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n244), .A3(new_n252), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n258), .B1(new_n267), .B2(new_n217), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n255), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n263), .B(KEYINPUT32), .C1(new_n269), .C2(new_n202), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT33), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n269), .B2(new_n202), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT71), .ZN(new_n274));
  XOR2_X1   g073(.A(G71gat), .B(G99gat), .Z(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n262), .A2(new_n270), .A3(new_n272), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n260), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n276), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n270), .A4(new_n262), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(KEYINPUT32), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n276), .A2(new_n271), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n202), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT34), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT36), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n294), .A3(new_n288), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n294), .B1(new_n284), .B2(new_n288), .ZN(new_n299));
  AOI211_X1 g098(.A(new_n291), .B(new_n287), .C1(new_n280), .C2(new_n283), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n210), .A2(new_n212), .B1(new_n215), .B2(new_n211), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n305), .B1(KEYINPUT2), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT2), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n304), .B2(KEYINPUT78), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n318), .A3(new_n309), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n303), .B(new_n311), .C1(new_n315), .C2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n311), .B1(new_n320), .B2(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n217), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT79), .Z(new_n326));
  AOI21_X1  g125(.A(new_n302), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n303), .B1(new_n322), .B2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n331), .B(new_n311), .C1(new_n320), .C2(new_n315), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n311), .C1(new_n320), .C2(new_n315), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n303), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n328), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n327), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n217), .A2(new_n322), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n330), .A2(new_n332), .B1(new_n341), .B2(KEYINPUT4), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n328), .ZN(new_n343));
  INV_X1    g142(.A(new_n326), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n302), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n340), .A2(new_n345), .A3(new_n350), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n352), .A2(KEYINPUT81), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n346), .B(new_n351), .C1(new_n356), .C2(KEYINPUT6), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT22), .ZN(new_n360));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n361), .B(new_n359), .C1(KEYINPUT22), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n266), .A2(new_n244), .A3(new_n252), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n265), .A2(new_n252), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(KEYINPUT29), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n368), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n375), .B1(new_n253), .B2(new_n254), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n371), .ZN(new_n380));
  INV_X1    g179(.A(new_n368), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n378), .A2(new_n382), .A3(new_n390), .A4(new_n386), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n385), .B(KEYINPUT74), .Z(new_n393));
  OR2_X1    g192(.A1(new_n374), .A2(new_n376), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n381), .B1(new_n394), .B2(new_n372), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n379), .A2(new_n381), .A3(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT75), .B(new_n393), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n387), .A2(new_n389), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n358), .A2(new_n392), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(KEYINPUT31), .B(G50gat), .Z(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n368), .B1(new_n332), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n322), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT3), .B1(new_n368), .B2(new_n405), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n363), .B1(new_n367), .B2(KEYINPUT82), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n367), .A2(KEYINPUT82), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n331), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n335), .A2(new_n337), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n411), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G22gat), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n411), .B(new_n420), .C1(new_n417), .C2(new_n408), .ZN(new_n421));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n419), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n404), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(new_n404), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n403), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n296), .A2(new_n301), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n296), .A2(new_n301), .A3(new_n434), .A4(new_n431), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT40), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n344), .B1(new_n342), .B2(new_n343), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT39), .B1(new_n324), .B2(new_n326), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n350), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT39), .B(new_n344), .C1(new_n342), .C2(new_n343), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT84), .B(new_n436), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n438), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n342), .A2(new_n343), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n344), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT39), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n350), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n447), .A3(new_n352), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n350), .A3(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT84), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n426), .A2(new_n429), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n354), .A2(new_n353), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n352), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n346), .A2(new_n353), .A3(new_n351), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n388), .A2(new_n391), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n378), .A2(new_n382), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n385), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n378), .B2(new_n382), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT38), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n381), .B1(new_n373), .B2(new_n377), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n379), .A2(new_n380), .A3(new_n368), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(KEYINPUT37), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n461), .A2(new_n467), .A3(new_n468), .A4(new_n393), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n458), .A2(new_n459), .A3(new_n464), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n433), .A2(new_n435), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n403), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n292), .A2(new_n473), .A3(new_n295), .A4(new_n454), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n299), .A2(new_n300), .A3(new_n430), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT85), .B(KEYINPUT35), .Z(new_n476));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n457), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n452), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(KEYINPUT35), .A2(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT90), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G1gat), .ZN(new_n484));
  INV_X1    g283(.A(G1gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT21), .ZN(new_n489));
  XOR2_X1   g288(.A(G71gat), .B(G78gat), .Z(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT94), .ZN(new_n491));
  XNOR2_X1  g290(.A(G71gat), .B(G78gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G57gat), .ZN(new_n497));
  OR2_X1    g296(.A1(KEYINPUT92), .A2(G64gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT92), .A2(G64gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT93), .B1(new_n497), .B2(G64gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G57gat), .B(G64gat), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT9), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n490), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n488), .B1(new_n489), .B2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT95), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n513));
  INV_X1    g312(.A(G231gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n509), .B(new_n489), .C1(new_n514), .C2(new_n370), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n370), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n496), .A2(new_n504), .B1(new_n490), .B2(new_n507), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(KEYINPUT21), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n521), .A2(new_n522), .A3(new_n513), .ZN(new_n525));
  XOR2_X1   g324(.A(G183gat), .B(G211gat), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n525), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n529), .B2(new_n523), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n512), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n523), .A3(new_n526), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n511), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n544), .A2(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT87), .ZN(new_n553));
  OR2_X1    g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(KEYINPUT14), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  XOR2_X1   g355(.A(G43gat), .B(G50gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n555), .A2(KEYINPUT15), .A3(new_n556), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n557), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n551), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n565), .A2(new_n551), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n536), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n571), .A2(new_n574), .A3(new_n536), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT97), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n571), .ZN(new_n579));
  INV_X1    g378(.A(new_n536), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n575), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  OAI211_X1 g387(.A(KEYINPUT97), .B(new_n588), .C1(new_n576), .C2(new_n577), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n535), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n517), .A2(new_n546), .A3(new_n549), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n595), .B(new_n596), .C1(new_n551), .C2(new_n517), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n551), .A2(KEYINPUT10), .A3(new_n517), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n594), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n595), .B1(new_n551), .B2(new_n517), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n594), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n592), .B1(new_n603), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n597), .A2(new_n601), .A3(new_n598), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n601), .B1(new_n597), .B2(new_n598), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n593), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT99), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n609), .B1(new_n619), .B2(new_n605), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n623), .B(new_n620), .C1(new_n611), .C2(new_n616), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G113gat), .B(G141gat), .Z(new_n627));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n488), .A2(new_n568), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n566), .A2(new_n570), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n488), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT91), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(KEYINPUT18), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n488), .B(new_n568), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n637), .B(KEYINPUT13), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT18), .B1(new_n635), .B2(new_n637), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n632), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n635), .A2(new_n637), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n632), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n647), .A2(new_n638), .A3(new_n641), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n481), .A2(new_n591), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n358), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n485), .ZN(G1324gat));
  INV_X1    g454(.A(new_n452), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g460(.A(KEYINPUT42), .B(new_n659), .S(new_n661), .Z(G1325gat));
  NAND2_X1  g461(.A1(new_n296), .A2(new_n301), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n299), .A2(new_n300), .ZN(new_n666));
  INV_X1    g465(.A(G15gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n653), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n454), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(new_n590), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n472), .B2(new_n480), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n531), .A2(new_n534), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(new_n626), .A3(new_n651), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n358), .A2(G29gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT101), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n481), .B2(new_n590), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n431), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n403), .A2(new_n430), .A3(KEYINPUT102), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n689), .A2(new_n471), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n691), .A2(new_n296), .A3(new_n301), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n686), .B(new_n590), .C1(new_n479), .C2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n296), .A3(new_n301), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n697));
  INV_X1    g496(.A(new_n478), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n299), .A2(new_n300), .A3(new_n430), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n700), .A2(KEYINPUT103), .A3(new_n686), .A4(new_n590), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n687), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n358), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n676), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G29gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n682), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n685), .A2(new_n706), .A3(new_n707), .ZN(G1328gat));
  OAI211_X1 g507(.A(new_n452), .B(new_n676), .C1(new_n687), .C2(new_n702), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G36gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n656), .A2(G36gat), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n481), .A2(new_n590), .A3(new_n676), .A4(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n674), .A2(KEYINPUT104), .A3(new_n676), .A4(new_n711), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT46), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n710), .B(KEYINPUT105), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n664), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n676), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n674), .A2(new_n666), .A3(new_n676), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n727), .A2(new_n723), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n725), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n454), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n703), .A2(new_n676), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n677), .A2(new_n430), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n732), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n737));
  AND3_X1   g536(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n734), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1331gat));
  NAND3_X1  g539(.A1(new_n675), .A2(new_n673), .A3(new_n651), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n625), .B(new_n741), .C1(new_n480), .C2(new_n696), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n704), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g543(.A(new_n452), .B(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n748), .B2(new_n747), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n742), .A2(G71gat), .A3(new_n663), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n742), .A2(new_n666), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(G71gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n742), .A2(new_n430), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n535), .A2(new_n651), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT109), .Z(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(new_n626), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n703), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n358), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n700), .A2(new_n590), .A3(new_n759), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n626), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n704), .A2(new_n538), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  OAI211_X1 g567(.A(new_n452), .B(new_n760), .C1(new_n687), .C2(new_n702), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G92gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n746), .A2(new_n539), .A3(new_n626), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n746), .B(new_n760), .C1(new_n687), .C2(new_n702), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n765), .B2(new_n772), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n777), .A2(KEYINPUT111), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  XNOR2_X1  g580(.A(KEYINPUT112), .B(G99gat), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n666), .A3(new_n626), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n761), .A2(new_n664), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(G1338gat));
  OAI211_X1 g584(.A(new_n430), .B(new_n760), .C1(new_n687), .C2(new_n702), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n454), .A2(G106gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n765), .A2(new_n626), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n787), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n741), .A2(new_n626), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n609), .B1(new_n618), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT54), .B1(new_n599), .B2(new_n593), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n603), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT114), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n614), .B(KEYINPUT54), .C1(new_n593), .C2(new_n599), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT55), .A4(new_n797), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n800), .A2(new_n799), .B1(new_n611), .B2(new_n616), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(new_n650), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n631), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n635), .A2(new_n637), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n639), .A2(new_n640), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n649), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n603), .A2(new_n592), .A3(new_n610), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT99), .B1(new_n614), .B2(new_n615), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n621), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n623), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n617), .A2(KEYINPUT100), .A3(new_n621), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n673), .B1(new_n807), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n649), .A2(new_n811), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n590), .A2(new_n820), .A3(new_n805), .A4(new_n806), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n622), .B2(new_n624), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n650), .A3(new_n806), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n590), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n590), .A2(new_n805), .A3(new_n820), .A4(new_n806), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT115), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n795), .B1(new_n829), .B2(new_n535), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n358), .A3(new_n746), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n475), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(new_n203), .A3(new_n651), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n830), .A2(new_n358), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n475), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n675), .B1(new_n823), .B2(new_n828), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n704), .B(new_n475), .C1(new_n837), .C2(new_n795), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n746), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n650), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n833), .B1(new_n841), .B2(new_n203), .ZN(G1340gat));
  NAND2_X1  g641(.A1(new_n626), .A2(new_n206), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G120gat), .B1(new_n832), .B2(new_n625), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(new_n832), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(G127gat), .A3(new_n675), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n840), .A2(new_n675), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  AOI21_X1  g650(.A(G127gat), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n840), .A2(new_n675), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n852), .B2(new_n854), .ZN(G1342gat));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n839), .ZN(new_n856));
  INV_X1    g655(.A(G134gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n590), .A2(new_n656), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT119), .Z(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n832), .B2(new_n673), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n861), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n861), .B2(KEYINPUT56), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n663), .A2(new_n358), .A3(new_n746), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n430), .B1(new_n837), .B2(new_n795), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(KEYINPUT121), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n675), .B1(new_n819), .B2(new_n821), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT57), .B(new_n430), .C1(new_n871), .C2(new_n795), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT121), .B1(new_n868), .B2(new_n869), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n650), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G141gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n663), .A2(new_n454), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n831), .A2(new_n306), .A3(new_n650), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1344gat));
  NOR2_X1   g682(.A1(new_n307), .A2(KEYINPUT59), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n625), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n430), .A2(new_n869), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n741), .B2(new_n626), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n591), .A2(KEYINPUT122), .A3(new_n625), .A4(new_n651), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n871), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(new_n626), .A3(new_n867), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT59), .B1(new_n895), .B2(new_n307), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n834), .A2(new_n877), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(new_n307), .A3(new_n626), .A4(new_n745), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1345gat));
  OR3_X1    g699(.A1(new_n885), .A2(new_n312), .A3(new_n535), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n831), .A2(new_n675), .A3(new_n877), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n312), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n885), .B2(new_n673), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n313), .A3(new_n860), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  INV_X1    g706(.A(new_n830), .ZN(new_n908));
  INV_X1    g707(.A(new_n475), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n704), .A3(new_n656), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n908), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G169gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n651), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n830), .A2(new_n704), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n475), .A2(new_n746), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n650), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n917), .A2(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n915), .B2(new_n625), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n625), .A2(G176gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n921), .B2(new_n926), .ZN(G1349gat));
  OAI21_X1  g726(.A(G183gat), .B1(new_n915), .B2(new_n535), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n922), .A2(new_n248), .A3(new_n675), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n249), .A3(new_n590), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n913), .A2(new_n590), .A3(new_n914), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n936), .A2(new_n937), .A3(G190gat), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n936), .B2(G190gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n663), .A2(new_n454), .A3(new_n745), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n918), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n650), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n663), .A2(new_n704), .A3(new_n656), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n894), .B2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n946), .B(new_n893), .C1(new_n868), .C2(KEYINPUT57), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n650), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  XOR2_X1   g749(.A(KEYINPUT126), .B(G204gat), .Z(new_n951));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n626), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NOR3_X1   g752(.A1(new_n945), .A2(new_n947), .A3(new_n625), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n951), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n894), .A2(new_n675), .A3(new_n944), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G211gat), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n364), .A3(new_n675), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1354gat));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n945), .B2(new_n947), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n590), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT127), .ZN(new_n963));
  OAI21_X1  g762(.A(G218gat), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n942), .A2(new_n365), .A3(new_n590), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


