//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT5), .ZN(new_n245));
  OAI21_X1  g0045(.A(KEYINPUT80), .B1(new_n245), .B2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT80), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n203), .B(G45), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n253), .C2(new_n248), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n250), .A2(new_n252), .A3(G274), .A4(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n245), .A2(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n254), .B(G270), .C1(new_n251), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT74), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT74), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n258), .A3(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G257), .A2(G1698), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n218), .B2(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n263), .A2(new_n265), .B1(G303), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n255), .B(new_n257), .C1(new_n269), .C2(new_n254), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G169), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT21), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n270), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n210), .ZN(new_n276));
  INV_X1    g0076(.A(G116), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G283), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n204), .C1(G33), .C2(new_n223), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT20), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(KEYINPUT20), .A3(new_n281), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT82), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(KEYINPUT82), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n275), .A2(new_n210), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n277), .B1(new_n203), .B2(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G116), .B2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n274), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n286), .B2(new_n287), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n270), .A2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n303), .B(new_n304), .C1(new_n270), .C2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n272), .B1(new_n303), .B2(new_n271), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n302), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n254), .A2(new_n314), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(G226), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT3), .B(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G222), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G223), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n312), .C1(G77), .C2(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT65), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n318), .A2(KEYINPUT65), .A3(new_n324), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n293), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n276), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n204), .A2(G1), .ZN(new_n334));
  INV_X1    g0134(.A(G50), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n333), .A2(new_n336), .B1(new_n335), .B2(new_n332), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G50), .A2(G58), .ZN(new_n338));
  INV_X1    g0138(.A(G68), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n204), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n204), .A2(new_n253), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n221), .A2(KEYINPUT8), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n221), .A2(KEYINPUT8), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n204), .A2(G33), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n340), .B(new_n343), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n337), .B1(new_n349), .B2(new_n296), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n327), .A2(new_n328), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n273), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n331), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT68), .B(G200), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n327), .A2(new_n356), .A3(new_n328), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT70), .ZN(new_n358));
  OAI211_X1 g0158(.A(KEYINPUT9), .B(new_n337), .C1(new_n349), .C2(new_n296), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT69), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT70), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n327), .A2(new_n365), .A3(new_n356), .A4(new_n328), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n350), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n368), .C1(new_n329), .C2(new_n305), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT10), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(KEYINPUT70), .A2(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n351), .A2(G190), .B1(new_n367), .B2(new_n350), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n366), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n354), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n339), .A2(G20), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(new_n347), .B2(new_n215), .C1(new_n335), .C2(new_n341), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n276), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT11), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT72), .B(KEYINPUT12), .Z(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n295), .B2(G68), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n290), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n295), .A2(new_n296), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n385), .A2(KEYINPUT71), .A3(new_n339), .A4(new_n334), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  INV_X1    g0187(.A(new_n385), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n334), .A2(new_n339), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n379), .B(new_n384), .C1(new_n386), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n222), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n319), .B(new_n392), .C1(G226), .C2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n254), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n314), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n254), .A3(G274), .ZN(new_n398));
  INV_X1    g0198(.A(G238), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n316), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n395), .B2(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G169), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(G179), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n405), .B2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n405), .A2(new_n305), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n412), .A2(new_n391), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT73), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n319), .A2(G232), .A3(new_n321), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT66), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n268), .A2(new_n399), .A3(new_n321), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G107), .B2(new_n268), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n254), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n398), .B1(new_n316), .B2(new_n216), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n273), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n295), .A2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n348), .B1(G20), .B2(G77), .ZN(new_n431));
  INV_X1    g0231(.A(new_n346), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n341), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n433), .B2(new_n276), .ZN(new_n434));
  INV_X1    g0234(.A(new_n334), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n388), .A2(G77), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n330), .B1(new_n424), .B2(new_n425), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n427), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n356), .B1(new_n424), .B2(new_n425), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n426), .B2(G190), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n411), .A2(new_n416), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n375), .A2(new_n418), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n398), .B1(new_n316), .B2(new_n222), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  MUX2_X1   g0247(.A(G223), .B(G226), .S(G1698), .Z(new_n448));
  AOI22_X1  g0248(.A1(new_n263), .A2(new_n448), .B1(G33), .B2(G87), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n308), .C1(new_n254), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n254), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n446), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(G200), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n346), .A2(new_n435), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n333), .B1(new_n332), .B2(new_n432), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n221), .A2(new_n339), .ZN(new_n457));
  NOR2_X1   g0257(.A1(G58), .A2(G68), .ZN(new_n458));
  OAI21_X1  g0258(.A(G20), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n204), .A2(new_n253), .A3(G159), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n261), .B1(new_n258), .B2(G33), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n253), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n266), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT7), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n204), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT7), .B1(new_n263), .B2(G20), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(G68), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT75), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n469), .A2(new_n470), .A3(new_n473), .A4(G68), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n464), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n468), .A2(new_n204), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n319), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT76), .B1(new_n258), .B2(G33), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT76), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n253), .A3(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n480), .A3(new_n267), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n204), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(KEYINPUT7), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n461), .B1(new_n483), .B2(G68), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n276), .B1(new_n484), .B2(KEYINPUT16), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n453), .B(new_n456), .C1(new_n475), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT78), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT17), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n488), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n489), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n456), .B1(new_n475), .B2(new_n485), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT18), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n452), .A2(G179), .ZN(new_n496));
  OAI21_X1  g0296(.A(G169), .B1(new_n451), .B2(new_n446), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n495), .B1(new_n494), .B2(new_n498), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n445), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n293), .A2(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n203), .A2(G33), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n296), .A2(new_n293), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n508), .B2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n483), .A2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n512), .A2(new_n223), .A3(G107), .ZN(new_n513));
  XNOR2_X1  g0313(.A(G97), .B(G107), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n515), .A2(new_n204), .B1(new_n215), .B2(new_n341), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n510), .B1(new_n518), .B2(new_n276), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n321), .A2(G244), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n467), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n321), .A2(KEYINPUT4), .A3(G244), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n268), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n524), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n319), .A2(new_n526), .A3(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n266), .A2(new_n267), .A3(G250), .A4(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n280), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n522), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n312), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n254), .B(G257), .C1(new_n251), .C2(new_n256), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n255), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(G200), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n530), .B1(new_n525), .B2(new_n527), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n254), .B1(new_n538), .B2(new_n522), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(G190), .A3(new_n535), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n519), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n542));
  OR2_X1    g0342(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n204), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n217), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n253), .A2(new_n277), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n204), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G20), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT22), .B1(new_n319), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n260), .A2(new_n262), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(KEYINPUT22), .A3(new_n266), .A4(new_n552), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n543), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  INV_X1    g0358(.A(new_n552), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n268), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n545), .A2(new_n546), .B1(new_n548), .B2(new_n204), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n543), .A2(new_n556), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n542), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n276), .ZN(new_n564));
  OR3_X1    g0364(.A1(new_n293), .A2(KEYINPUT84), .A3(G107), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT84), .B1(new_n293), .B2(G107), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(G107), .B2(new_n508), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G250), .A2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n224), .B2(G1698), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n263), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n253), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n312), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n254), .B(G264), .C1(new_n251), .C2(new_n256), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(new_n305), .A3(new_n255), .A4(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n263), .A2(new_n572), .B1(G33), .B2(G294), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n255), .B(new_n577), .C1(new_n579), .C2(new_n254), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n413), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n564), .A2(new_n570), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n516), .B1(G107), .B2(new_n483), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n509), .B1(new_n584), .B2(new_n296), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n533), .A2(new_n273), .A3(new_n536), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n330), .B1(new_n539), .B2(new_n535), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n541), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n330), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G179), .B2(new_n580), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n564), .B2(new_n570), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n203), .A2(new_n313), .A3(G45), .ZN(new_n593));
  INV_X1    g0393(.A(G45), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(G1), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n254), .B(new_n593), .C1(G250), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G238), .A2(G1698), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n216), .B2(G1698), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n548), .B1(new_n263), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n254), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n355), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n305), .B(new_n596), .C1(new_n599), .C2(new_n254), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n394), .B2(new_n204), .ZN(new_n605));
  NOR4_X1   g0405(.A1(KEYINPUT81), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT81), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G87), .A2(G97), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n217), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n339), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n555), .A2(new_n266), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n604), .B1(new_n347), .B2(new_n223), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n276), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n508), .A2(G87), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n295), .A2(new_n430), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n603), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n600), .A2(new_n330), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n273), .B(new_n596), .C1(new_n599), .C2(new_n254), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n618), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n507), .A2(new_n429), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n592), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n311), .A2(new_n504), .A3(new_n589), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n439), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n411), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n493), .A2(new_n416), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n502), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n370), .A2(new_n374), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n354), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n504), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .A3(new_n620), .A4(new_n625), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n615), .A2(KEYINPUT85), .A3(new_n616), .A4(new_n618), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n640), .A2(new_n641), .B1(new_n601), .B2(new_n602), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n621), .A2(new_n622), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n617), .B(new_n624), .C1(new_n614), .C2(new_n276), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n642), .A2(new_n588), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n637), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n302), .A2(new_n310), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n592), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n641), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n650), .B2(new_n603), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n588), .A3(new_n541), .A4(new_n583), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n647), .B(new_n625), .C1(new_n649), .C2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n634), .B1(new_n635), .B2(new_n654), .ZN(G369));
  NAND2_X1  g0455(.A1(new_n290), .A2(new_n204), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n311), .B1(new_n303), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n648), .A2(new_n301), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n592), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n564), .A2(new_n570), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n668), .A3(new_n583), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n666), .B2(new_n662), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(G330), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n648), .A2(new_n662), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n592), .A2(new_n662), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n207), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n606), .A2(new_n609), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n277), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n203), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n213), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT88), .Z(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n589), .A2(new_n311), .A3(new_n627), .A4(new_n662), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n535), .B1(new_n532), .B2(new_n312), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n577), .B1(new_n579), .B2(new_n254), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n600), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n263), .A2(new_n265), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n268), .A2(G303), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n254), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n255), .A2(new_n257), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n273), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n533), .A2(new_n536), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n600), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT89), .B(new_n596), .C1(new_n599), .C2(new_n254), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n270), .A2(new_n273), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n701), .A2(new_n705), .A3(new_n706), .A4(new_n580), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n690), .A2(new_n692), .A3(new_n697), .A4(KEYINPUT30), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n700), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n661), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n689), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n653), .A2(new_n662), .ZN(new_n717));
  XNOR2_X1  g0517(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n541), .A2(new_n583), .A3(new_n588), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n650), .A2(new_n603), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n625), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n666), .A2(new_n302), .A3(new_n310), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n645), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT26), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n626), .B2(new_n588), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT91), .B(new_n726), .C1(new_n626), .C2(new_n588), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n651), .A2(new_n636), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n729), .B(new_n730), .C1(new_n726), .C2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n661), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n716), .B1(new_n719), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n688), .B1(new_n735), .B2(G1), .ZN(G364));
  NAND2_X1  g0536(.A1(new_n665), .A2(G330), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n289), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n203), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n738), .B1(G330), .B2(new_n665), .C1(new_n681), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(new_n741), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n680), .A2(new_n268), .ZN(new_n744));
  NAND2_X1  g0544(.A1(G355), .A2(KEYINPUT93), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G355), .A2(KEYINPUT93), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n207), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n680), .A2(new_n263), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n594), .B2(new_n685), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n240), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n210), .B1(G20), .B2(new_n330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  OAI21_X1  g0559(.A(new_n743), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n355), .A2(new_n204), .A3(G179), .A4(new_n305), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n268), .B1(new_n761), .B2(G87), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n204), .B1(new_n765), .B2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n223), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n204), .A2(new_n273), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n413), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n771), .A2(new_n215), .B1(new_n774), .B2(new_n339), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n308), .A2(new_n772), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n767), .B(new_n775), .C1(G50), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n204), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n765), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n356), .A2(new_n273), .A3(new_n778), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G107), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n777), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n308), .A2(new_n769), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT95), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT95), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n764), .B(new_n786), .C1(G58), .C2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n761), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n783), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n319), .B1(new_n799), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n771), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  OAI22_X1  g0603(.A1(new_n774), .A2(new_n803), .B1(new_n574), .B2(new_n766), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n798), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  INV_X1    g0606(.A(G326), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n776), .B(KEYINPUT98), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n805), .B1(new_n806), .B2(new_n790), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n793), .A2(new_n794), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n760), .B1(new_n810), .B2(new_n757), .ZN(new_n811));
  INV_X1    g0611(.A(new_n756), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n665), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n742), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  INV_X1    g0615(.A(new_n757), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n755), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n784), .A2(G87), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n319), .B1(new_n799), .B2(G311), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n223), .C2(new_n766), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n776), .A2(G303), .B1(new_n770), .B2(G116), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n797), .B2(new_n774), .C1(new_n790), .C2(new_n574), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G107), .C2(new_n761), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n776), .A2(G137), .B1(new_n773), .B2(G150), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n780), .B2(new_n771), .C1(new_n790), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n263), .B1(new_n221), .B2(new_n766), .C1(new_n828), .C2(new_n779), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n783), .A2(new_n339), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(G50), .C2(new_n761), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n823), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n743), .B1(G77), .B2(new_n817), .C1(new_n832), .C2(new_n816), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  NAND4_X1  g0634(.A1(new_n662), .A2(new_n427), .A3(new_n437), .A4(new_n438), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n441), .A2(new_n440), .B1(new_n437), .B2(new_n661), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n439), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n834), .B1(new_n754), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n441), .A2(new_n440), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n839), .A2(new_n439), .A3(new_n661), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n625), .B1(new_n652), .B2(new_n649), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n626), .A2(new_n588), .A3(new_n726), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n731), .B2(new_n726), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n717), .ZN(new_n845));
  INV_X1    g0645(.A(new_n837), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(new_n715), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n743), .B1(new_n847), .B2(new_n715), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n739), .A2(new_n203), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n719), .A2(new_n734), .A3(new_n504), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n634), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT103), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n494), .A2(new_n498), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n494), .A2(new_n659), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n486), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n467), .A2(new_n204), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n339), .B1(new_n862), .B2(KEYINPUT7), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n473), .B1(new_n863), .B2(new_n469), .ZN(new_n864));
  INV_X1    g0664(.A(new_n474), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n463), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n276), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n472), .A2(new_n474), .ZN(new_n868));
  INV_X1    g0668(.A(new_n461), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n456), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n659), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n498), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n486), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n861), .B1(new_n874), .B2(KEYINPUT37), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n493), .B2(new_n502), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n857), .A2(new_n486), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n879), .A2(KEYINPUT102), .A3(new_n859), .A4(new_n858), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n860), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n456), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n482), .A2(KEYINPUT7), .ZN(new_n884));
  INV_X1    g0684(.A(new_n477), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(G68), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n869), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n296), .B1(new_n887), .B2(new_n462), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n883), .B1(new_n866), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n498), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n486), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n659), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n880), .A2(new_n882), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n490), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n489), .B1(new_n486), .B2(new_n491), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n857), .A2(KEYINPUT18), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n499), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n893), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n856), .B1(new_n878), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n405), .A2(G169), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT14), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n408), .A3(new_n407), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n391), .A3(new_n662), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n909));
  INV_X1    g0709(.A(new_n872), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n898), .B2(new_n900), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n871), .A2(new_n498), .B1(new_n889), .B2(new_n453), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n859), .B1(new_n912), .B2(new_n872), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n911), .B(KEYINPUT38), .C1(new_n913), .C2(new_n861), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n903), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n909), .A2(new_n914), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n661), .A2(new_n391), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n411), .A2(new_n416), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n391), .B(new_n661), .C1(new_n906), .C2(new_n415), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n835), .B(KEYINPUT101), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n844), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n917), .A2(new_n925), .B1(new_n900), .B2(new_n892), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n855), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(G330), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n909), .A2(new_n914), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n709), .A2(new_n933), .A3(KEYINPUT31), .A4(new_n661), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n689), .A2(new_n932), .A3(new_n712), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n837), .B1(new_n919), .B2(new_n920), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT40), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n878), .B2(new_n902), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n935), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n635), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n929), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n852), .B1(new_n928), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n928), .B2(new_n949), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT35), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n515), .A2(new_n952), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n277), .B(new_n212), .C1(new_n515), .C2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n953), .B1(new_n955), .B2(KEYINPUT100), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT100), .B2(new_n955), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n457), .A2(new_n213), .A3(new_n215), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n339), .A2(G50), .ZN(new_n960));
  OAI211_X1 g0760(.A(G1), .B(new_n289), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n951), .A2(new_n958), .A3(new_n961), .ZN(G367));
  NAND3_X1  g0762(.A1(new_n661), .A2(new_n640), .A3(new_n641), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(new_n625), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n651), .A2(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n756), .ZN(new_n970));
  INV_X1    g0770(.A(new_n759), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n207), .B2(new_n429), .C1(new_n236), .C2(new_n750), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n743), .ZN(new_n973));
  INV_X1    g0773(.A(G137), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n319), .B1(new_n974), .B2(new_n779), .C1(new_n774), .C2(new_n780), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n795), .A2(new_n221), .B1(new_n215), .B2(new_n783), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n771), .A2(new_n335), .B1(new_n766), .B2(new_n339), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n825), .B2(new_n808), .C1(new_n342), .C2(new_n790), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT46), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n761), .A2(G116), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n791), .A2(G303), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n980), .B2(new_n981), .C1(new_n801), .C2(new_n808), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n784), .A2(G97), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G283), .A2(new_n770), .B1(new_n773), .B2(G294), .ZN(new_n985));
  INV_X1    g0785(.A(new_n766), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(G107), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n263), .B1(G317), .B2(new_n799), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n979), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n973), .B1(new_n992), .B2(new_n757), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n970), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n541), .B(new_n588), .C1(new_n662), .C2(new_n519), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n636), .A2(new_n661), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n677), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n677), .A2(new_n998), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n672), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n672), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n674), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n675), .B1(new_n670), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n737), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n738), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n735), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n735), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n681), .B(KEYINPUT41), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n741), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n673), .A2(new_n998), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n675), .A2(new_n998), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT107), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1018), .B2(KEYINPUT42), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n995), .A2(new_n666), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n661), .B1(new_n1023), .B2(new_n588), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1018), .B2(KEYINPUT42), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1022), .A2(new_n1025), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT43), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n969), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1022), .A2(new_n1027), .A3(new_n969), .A4(new_n1025), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n1017), .A3(new_n1030), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1016), .A2(new_n1034), .A3(KEYINPUT108), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n735), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1006), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n1004), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1039), .B2(new_n1011), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n740), .B1(new_n1040), .B2(new_n1014), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1033), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n1031), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1036), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n994), .B1(new_n1035), .B2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n1011), .A2(new_n741), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1011), .A2(new_n735), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1012), .A2(new_n681), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n233), .A2(new_n594), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(new_n749), .B1(new_n683), .B2(new_n744), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n346), .A2(new_n335), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n594), .B1(new_n339), .B2(new_n215), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1052), .A2(new_n683), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1050), .A2(new_n1054), .B1(G107), .B2(new_n207), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n971), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G68), .A2(new_n770), .B1(new_n773), .B2(new_n346), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n986), .A2(new_n430), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n776), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1058), .C1(new_n780), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n467), .B1(G150), .B2(new_n799), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n984), .B(new_n1061), .C1(new_n215), .C2(new_n795), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(G50), .C2(new_n791), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n761), .A2(G294), .B1(G283), .B2(new_n986), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G303), .A2(new_n770), .B1(new_n773), .B2(G311), .ZN(new_n1065));
  INV_X1    g0865(.A(G317), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n808), .B2(new_n806), .C1(new_n1066), .C2(new_n790), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT110), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n467), .B1(new_n807), .B2(new_n779), .C1(new_n783), .C2(new_n277), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT111), .Z(new_n1075));
  AOI21_X1  g0875(.A(new_n1063), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n743), .B(new_n1056), .C1(new_n1076), .C2(new_n816), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT112), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n670), .B2(new_n812), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .C1(new_n1080), .C2(new_n1081), .ZN(G393));
  NAND3_X1  g0882(.A1(new_n1039), .A2(new_n735), .A3(new_n1011), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n681), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n998), .A2(new_n756), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n971), .B1(new_n223), .B2(new_n207), .C1(new_n243), .C2(new_n750), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(KEYINPUT113), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT113), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n743), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n790), .A2(new_n801), .B1(new_n1066), .B2(new_n1059), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT52), .Z(new_n1092));
  OAI221_X1 g0892(.A(new_n268), .B1(new_n806), .B2(new_n779), .C1(new_n774), .C2(new_n796), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n771), .A2(new_n574), .B1(new_n766), .B2(new_n277), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n785), .B1(new_n797), .B2(new_n795), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n790), .A2(new_n780), .B1(new_n342), .B2(new_n1059), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  AOI22_X1  g0898(.A1(G50), .A2(new_n773), .B1(new_n770), .B2(new_n346), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n215), .B2(new_n766), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT114), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n467), .B1(G143), .B2(new_n799), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n818), .B(new_n1102), .C1(new_n339), .C2(new_n795), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1098), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1088), .B(new_n1090), .C1(new_n1105), .C2(new_n757), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1039), .A2(new_n741), .B1(new_n1086), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1107), .ZN(G390));
  INV_X1    g0908(.A(new_n681), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n894), .B1(new_n881), .B2(new_n860), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n882), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n901), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n877), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n914), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n836), .A2(new_n439), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n733), .A2(new_n1116), .B1(new_n439), .B2(new_n662), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1114), .B(new_n907), .C1(new_n1117), .C2(new_n922), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n714), .A2(G330), .A3(new_n846), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n921), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT39), .B1(new_n1113), .B2(new_n914), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n925), .B2(new_n908), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n923), .B1(new_n653), .B2(new_n840), .ZN(new_n1127));
  OAI211_X1 g0927(.A(KEYINPUT115), .B(new_n907), .C1(new_n1127), .C2(new_n922), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1118), .B(new_n1121), .C1(new_n1124), .C2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n903), .A2(new_n915), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n733), .A2(new_n1116), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n835), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n908), .B1(new_n1134), .B2(new_n921), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1131), .A2(new_n1132), .B1(new_n1135), .B2(new_n1114), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n935), .A2(new_n936), .A3(G330), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n946), .A2(new_n929), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n504), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n853), .A2(new_n634), .A3(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n946), .A2(new_n929), .A3(new_n837), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1121), .B(new_n1117), .C1(new_n921), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1137), .B1(new_n1120), .B2(new_n921), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1127), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1141), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1109), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1130), .B(new_n1147), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n743), .B1(new_n346), .B2(new_n817), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n791), .A2(G116), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n830), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1059), .A2(new_n797), .B1(new_n771), .B2(new_n223), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G107), .B2(new_n773), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n268), .B1(new_n766), .B2(new_n215), .C1(new_n574), .C2(new_n779), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G87), .B2(new_n761), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1059), .A2(new_n1160), .B1(new_n780), .B2(new_n766), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G137), .B2(new_n773), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n268), .B1(new_n799), .B2(G125), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n771), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G50), .B2(new_n784), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1162), .B(new_n1166), .C1(new_n828), .C2(new_n790), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n761), .A2(G150), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1159), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1170), .B2(new_n757), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1124), .B2(new_n755), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1138), .B2(new_n740), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1151), .A2(new_n1173), .ZN(G378));
  INV_X1    g0974(.A(new_n1141), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1150), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n927), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n940), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT105), .B1(new_n935), .B2(new_n936), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT40), .B1(new_n1180), .B2(new_n917), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n944), .A2(G330), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n375), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n350), .A2(new_n659), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1184), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(new_n1183), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1181), .A2(new_n1182), .A3(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n929), .B1(new_n1114), .B2(new_n943), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n942), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1177), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1193), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n942), .A2(new_n1196), .A3(new_n1195), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n927), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(KEYINPUT118), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT118), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n1177), .C1(new_n1194), .C2(new_n1197), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1176), .A2(new_n1202), .A3(KEYINPUT57), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1176), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n681), .B(new_n1205), .C1(new_n1207), .C2(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n741), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n743), .B1(G50), .B2(new_n817), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n761), .A2(G77), .B1(G283), .B2(new_n799), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n263), .A2(G41), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n221), .C2(new_n783), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT116), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n773), .A2(G97), .B1(G68), .B2(new_n986), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n429), .B2(new_n771), .C1(new_n277), .C2(new_n1059), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G107), .B2(new_n791), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT117), .Z(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G33), .A2(G41), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1212), .A2(G50), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n766), .A2(new_n342), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n771), .A2(new_n974), .B1(new_n774), .B2(new_n828), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(G125), .C2(new_n776), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n1160), .B2(new_n790), .C1(new_n795), .C2(new_n1164), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n799), .A2(G124), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1222), .B(new_n1229), .C1(new_n783), .C2(new_n780), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1227), .B2(KEYINPUT59), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1223), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1220), .A2(new_n1221), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1210), .B1(new_n1233), .B2(new_n757), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1193), .B2(new_n755), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1209), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1208), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n922), .A2(new_n754), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n743), .B1(G68), .B2(new_n817), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n791), .A2(G137), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n761), .A2(G159), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n263), .B1(new_n1160), .B2(new_n779), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n784), .B2(G58), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1059), .A2(new_n828), .B1(new_n774), .B2(new_n1164), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n771), .A2(new_n342), .B1(new_n766), .B2(new_n335), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n791), .A2(G283), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n761), .A2(G97), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1059), .A2(new_n574), .B1(new_n771), .B2(new_n217), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G116), .B2(new_n773), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1058), .B(new_n268), .C1(new_n796), .C2(new_n779), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G77), .B2(new_n784), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1248), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1240), .B1(new_n1256), .B2(new_n757), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1238), .A2(new_n741), .B1(new_n1239), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1148), .A2(new_n1015), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1238), .A2(new_n1175), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT119), .Z(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G381));
  INV_X1    g1063(.A(new_n994), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT108), .B1(new_n1016), .B2(new_n1034), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1041), .A2(new_n1043), .A3(new_n1036), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(G390), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(G378), .A3(G375), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT120), .Z(G407));
  NOR2_X1   g1071(.A1(new_n1151), .A2(new_n1173), .ZN(new_n1272));
  INV_X1    g1072(.A(G343), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G375), .C2(new_n1274), .ZN(G409));
  XNOR2_X1  g1075(.A(G393), .B(new_n814), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n994), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1279), .B2(new_n1267), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(G390), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n994), .A3(new_n1277), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1276), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1280), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1273), .A2(G213), .A3(G2897), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1260), .B(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n681), .A3(new_n1148), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G384), .A3(new_n1258), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1291), .B2(new_n1258), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1292), .A3(new_n1287), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT122), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1202), .A2(new_n1204), .A3(new_n741), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1235), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1014), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT121), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1302), .A2(new_n1176), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1302), .B2(new_n1176), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1301), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1299), .B1(new_n1306), .B2(G378), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G378), .A2(new_n1208), .A3(new_n1236), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1305), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1302), .A2(new_n1176), .A3(new_n1303), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(KEYINPUT122), .B(new_n1272), .C1(new_n1311), .C2(new_n1301), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1307), .A2(new_n1308), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1273), .A2(G213), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1298), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1286), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  AOI211_X1 g1117(.A(KEYINPUT125), .B(new_n1298), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1320), .A4(new_n1314), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(KEYINPUT126), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1313), .A2(new_n1320), .A3(new_n1314), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT123), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT123), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1313), .A2(new_n1325), .A3(new_n1320), .A4(new_n1314), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1319), .A2(new_n1322), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT62), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1298), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1330), .B1(new_n1331), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1329), .A2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1272), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1308), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1340), .A2(new_n1320), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1320), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1330), .A3(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1343), .A2(KEYINPUT127), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(KEYINPUT127), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1330), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(G402));
endmodule


