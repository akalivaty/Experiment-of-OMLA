

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777;

  AND2_X1 U368 ( .A1(n640), .A2(n639), .ZN(n680) );
  NAND2_X1 U369 ( .A1(n359), .A2(n356), .ZN(n776) );
  XOR2_X1 U370 ( .A(KEYINPUT110), .B(n586), .Z(n733) );
  XNOR2_X1 U371 ( .A(n431), .B(n430), .ZN(n521) );
  AND2_X1 U372 ( .A1(n676), .A2(n465), .ZN(n431) );
  BUF_X1 U373 ( .A(G953), .Z(n345) );
  NOR2_X1 U374 ( .A1(n498), .A2(n416), .ZN(n417) );
  XNOR2_X1 U375 ( .A(G119), .B(G128), .ZN(n418) );
  BUF_X1 U376 ( .A(n453), .Z(n769) );
  INV_X1 U377 ( .A(G953), .ZN(n453) );
  XNOR2_X2 U378 ( .A(n601), .B(n353), .ZN(n735) );
  NAND2_X2 U379 ( .A1(n614), .A2(n735), .ZN(n582) );
  XNOR2_X2 U380 ( .A(n493), .B(n369), .ZN(n385) );
  NOR2_X2 U381 ( .A1(n653), .A2(n686), .ZN(n654) );
  NOR2_X2 U382 ( .A1(n646), .A2(n686), .ZN(n647) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n483) );
  XNOR2_X2 U384 ( .A(n469), .B(n468), .ZN(n604) );
  XNOR2_X2 U385 ( .A(n443), .B(n383), .ZN(n681) );
  XNOR2_X2 U386 ( .A(n455), .B(G134), .ZN(n493) );
  INV_X2 U387 ( .A(n560), .ZN(n775) );
  INV_X1 U388 ( .A(n482), .ZN(n369) );
  XNOR2_X1 U389 ( .A(n370), .B(KEYINPUT67), .ZN(n482) );
  INV_X1 U390 ( .A(G131), .ZN(n370) );
  AND2_X1 U391 ( .A1(n380), .A2(n379), .ZN(n663) );
  NAND2_X1 U392 ( .A1(n390), .A2(n388), .ZN(n387) );
  AND2_X1 U393 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U394 ( .A1(n538), .A2(n389), .ZN(n388) );
  AND2_X1 U395 ( .A1(n539), .A2(n566), .ZN(n389) );
  NOR2_X1 U396 ( .A1(n524), .A2(n688), .ZN(n531) );
  AND2_X1 U397 ( .A1(n393), .A2(n352), .ZN(n504) );
  XNOR2_X1 U398 ( .A(n550), .B(n549), .ZN(n777) );
  OR2_X2 U399 ( .A1(n374), .A2(n371), .ZN(n528) );
  NOR2_X1 U400 ( .A1(n508), .A2(n507), .ZN(n730) );
  XNOR2_X1 U401 ( .A(n434), .B(KEYINPUT75), .ZN(n506) );
  XNOR2_X1 U402 ( .A(n766), .B(KEYINPUT71), .ZN(n462) );
  XNOR2_X1 U403 ( .A(n451), .B(KEYINPUT69), .ZN(n384) );
  XNOR2_X1 U404 ( .A(n406), .B(n405), .ZN(n766) );
  XOR2_X1 U405 ( .A(KEYINPUT95), .B(G107), .Z(n405) );
  XNOR2_X1 U406 ( .A(G110), .B(G104), .ZN(n404) );
  XNOR2_X2 U407 ( .A(n582), .B(n581), .ZN(n629) );
  BUF_X1 U408 ( .A(n520), .Z(n346) );
  XNOR2_X1 U409 ( .A(KEYINPUT68), .B(G140), .ZN(n409) );
  AND2_X1 U410 ( .A1(n615), .A2(n655), .ZN(n616) );
  NAND2_X1 U411 ( .A1(n386), .A2(n365), .ZN(n596) );
  XOR2_X1 U412 ( .A(G140), .B(KEYINPUT12), .Z(n485) );
  XOR2_X1 U413 ( .A(G122), .B(G104), .Z(n480) );
  INV_X1 U414 ( .A(G146), .ZN(n413) );
  NAND2_X1 U415 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U416 ( .A1(n373), .A2(KEYINPUT0), .ZN(n372) );
  NAND2_X1 U417 ( .A1(n640), .A2(n348), .ZN(n381) );
  XNOR2_X1 U418 ( .A(n423), .B(n666), .ZN(n676) );
  INV_X1 U419 ( .A(KEYINPUT64), .ZN(n412) );
  INV_X1 U420 ( .A(G237), .ZN(n464) );
  NAND2_X1 U421 ( .A1(n476), .A2(n398), .ZN(n397) );
  NAND2_X1 U422 ( .A1(n604), .A2(n378), .ZN(n376) );
  NAND2_X1 U423 ( .A1(n475), .A2(n378), .ZN(n375) );
  XNOR2_X1 U424 ( .A(G116), .B(G107), .ZN(n494) );
  XNOR2_X1 U425 ( .A(G113), .B(G143), .ZN(n479) );
  XNOR2_X1 U426 ( .A(n411), .B(n462), .ZN(n383) );
  XNOR2_X1 U427 ( .A(n410), .B(n422), .ZN(n411) );
  XNOR2_X1 U428 ( .A(n377), .B(n519), .ZN(n548) );
  XNOR2_X1 U429 ( .A(n507), .B(n445), .ZN(n597) );
  AND2_X1 U430 ( .A1(n626), .A2(n382), .ZN(n628) );
  NAND2_X1 U431 ( .A1(n358), .A2(n593), .ZN(n357) );
  NOR2_X1 U432 ( .A1(n698), .A2(n583), .ZN(n364) );
  NOR2_X1 U433 ( .A1(n612), .A2(n382), .ZN(n613) );
  XNOR2_X1 U434 ( .A(n607), .B(n606), .ZN(n699) );
  INV_X1 U435 ( .A(KEYINPUT81), .ZN(n606) );
  XNOR2_X1 U436 ( .A(n381), .B(n661), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n368), .B(n676), .ZN(n367) );
  NAND2_X1 U438 ( .A1(n680), .A2(G217), .ZN(n368) );
  NAND2_X1 U439 ( .A1(n698), .A2(n583), .ZN(n347) );
  AND2_X1 U440 ( .A1(n639), .A2(G472), .ZN(n348) );
  XNOR2_X1 U441 ( .A(n525), .B(KEYINPUT1), .ZN(n520) );
  XOR2_X1 U442 ( .A(n440), .B(n439), .Z(n349) );
  AND2_X1 U443 ( .A1(n467), .A2(G210), .ZN(n350) );
  AND2_X1 U444 ( .A1(n605), .A2(n366), .ZN(n351) );
  AND2_X1 U445 ( .A1(n397), .A2(n400), .ZN(n352) );
  XOR2_X1 U446 ( .A(KEYINPUT74), .B(KEYINPUT38), .Z(n353) );
  INV_X1 U447 ( .A(KEYINPUT0), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n477), .B(KEYINPUT80), .ZN(n478) );
  AND2_X1 U449 ( .A1(n639), .A2(G210), .ZN(n354) );
  AND2_X1 U450 ( .A1(n639), .A2(G475), .ZN(n355) );
  NOR2_X1 U451 ( .A1(n769), .A2(G952), .ZN(n686) );
  INV_X1 U452 ( .A(n686), .ZN(n379) );
  OR2_X1 U453 ( .A1(n733), .A2(n357), .ZN(n356) );
  INV_X1 U454 ( .A(n605), .ZN(n358) );
  NOR2_X1 U455 ( .A1(n360), .A2(n351), .ZN(n359) );
  AND2_X1 U456 ( .A1(n733), .A2(n366), .ZN(n360) );
  NAND2_X1 U457 ( .A1(n362), .A2(n361), .ZN(n386) );
  NAND2_X1 U458 ( .A1(n629), .A2(KEYINPUT40), .ZN(n361) );
  NOR2_X1 U459 ( .A1(n363), .A2(n364), .ZN(n362) );
  NOR2_X1 U460 ( .A1(n629), .A2(n347), .ZN(n363) );
  INV_X1 U461 ( .A(n776), .ZN(n365) );
  INV_X1 U462 ( .A(n593), .ZN(n366) );
  AND2_X1 U463 ( .A1(n367), .A2(n379), .ZN(G66) );
  XNOR2_X2 U464 ( .A(G143), .B(G128), .ZN(n455) );
  NAND2_X2 U465 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X2 U466 ( .A1(n636), .A2(n637), .ZN(n640) );
  NOR2_X1 U467 ( .A1(n604), .A2(n372), .ZN(n371) );
  INV_X1 U468 ( .A(n475), .ZN(n373) );
  NAND2_X1 U469 ( .A1(n528), .A2(n516), .ZN(n377) );
  INV_X1 U470 ( .A(n601), .ZN(n382) );
  XNOR2_X2 U471 ( .A(n466), .B(n350), .ZN(n601) );
  XNOR2_X2 U472 ( .A(n667), .B(n413), .ZN(n443) );
  XNOR2_X2 U473 ( .A(n385), .B(n384), .ZN(n667) );
  NAND2_X1 U474 ( .A1(n640), .A2(n354), .ZN(n652) );
  NAND2_X1 U475 ( .A1(n640), .A2(n355), .ZN(n645) );
  XNOR2_X1 U476 ( .A(n386), .B(G131), .ZN(G33) );
  XNOR2_X2 U477 ( .A(n387), .B(n567), .ZN(n758) );
  NAND2_X1 U478 ( .A1(n558), .A2(n557), .ZN(n391) );
  NAND2_X1 U479 ( .A1(n562), .A2(n563), .ZN(n392) );
  NAND2_X1 U480 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U481 ( .A1(n717), .A2(n478), .ZN(n394) );
  NAND2_X1 U482 ( .A1(n396), .A2(n399), .ZN(n395) );
  INV_X1 U483 ( .A(n717), .ZN(n396) );
  XNOR2_X2 U484 ( .A(n448), .B(n447), .ZN(n717) );
  INV_X1 U485 ( .A(n478), .ZN(n398) );
  NAND2_X1 U486 ( .A1(n528), .A2(n478), .ZN(n399) );
  INV_X1 U487 ( .A(n612), .ZN(n400) );
  OR2_X1 U488 ( .A1(G902), .A2(n677), .ZN(n401) );
  XOR2_X1 U489 ( .A(G110), .B(KEYINPUT24), .Z(n402) );
  XOR2_X1 U490 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n403) );
  NAND2_X1 U491 ( .A1(n699), .A2(n608), .ZN(n611) );
  XNOR2_X1 U492 ( .A(n441), .B(n349), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n404), .B(G101), .ZN(n406) );
  XOR2_X1 U494 ( .A(KEYINPUT79), .B(KEYINPUT97), .Z(n408) );
  AND2_X1 U495 ( .A1(n769), .A2(G227), .ZN(n407) );
  XNOR2_X1 U496 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n409), .B(G137), .ZN(n422) );
  XNOR2_X1 U498 ( .A(n412), .B(KEYINPUT4), .ZN(n451) );
  OR2_X2 U499 ( .A1(n681), .A2(G902), .ZN(n414) );
  XNOR2_X2 U500 ( .A(n414), .B(G469), .ZN(n525) );
  NAND2_X1 U501 ( .A1(n453), .A2(G234), .ZN(n415) );
  XNOR2_X1 U502 ( .A(n415), .B(KEYINPUT8), .ZN(n498) );
  INV_X1 U503 ( .A(G221), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n417), .B(n402), .ZN(n420) );
  XNOR2_X1 U505 ( .A(n418), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U506 ( .A(n420), .B(n419), .ZN(n423) );
  XNOR2_X2 U507 ( .A(G146), .B(G125), .ZN(n450) );
  INV_X1 U508 ( .A(KEYINPUT10), .ZN(n421) );
  XNOR2_X1 U509 ( .A(n450), .B(n421), .ZN(n481) );
  XNOR2_X1 U510 ( .A(n481), .B(n422), .ZN(n666) );
  INV_X1 U511 ( .A(G902), .ZN(n465) );
  XNOR2_X1 U512 ( .A(KEYINPUT94), .B(KEYINPUT15), .ZN(n424) );
  XNOR2_X1 U513 ( .A(n424), .B(G902), .ZN(n638) );
  NAND2_X1 U514 ( .A1(n638), .A2(G234), .ZN(n425) );
  XNOR2_X1 U515 ( .A(KEYINPUT20), .B(n425), .ZN(n432) );
  NAND2_X1 U516 ( .A1(n432), .A2(G217), .ZN(n429) );
  XNOR2_X1 U517 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n427) );
  INV_X1 U518 ( .A(KEYINPUT25), .ZN(n426) );
  XNOR2_X1 U519 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U520 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U521 ( .A1(n432), .A2(G221), .ZN(n433) );
  XNOR2_X1 U522 ( .A(n433), .B(KEYINPUT21), .ZN(n721) );
  INV_X1 U523 ( .A(n721), .ZN(n588) );
  AND2_X1 U524 ( .A1(n521), .A2(n588), .ZN(n725) );
  NAND2_X1 U525 ( .A1(n520), .A2(n725), .ZN(n434) );
  INV_X1 U526 ( .A(KEYINPUT3), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n435), .B(G119), .ZN(n437) );
  XNOR2_X1 U528 ( .A(G116), .B(G113), .ZN(n436) );
  XNOR2_X1 U529 ( .A(n437), .B(n436), .ZN(n460) );
  NAND2_X1 U530 ( .A1(n483), .A2(G210), .ZN(n438) );
  XNOR2_X1 U531 ( .A(n460), .B(n438), .ZN(n441) );
  XOR2_X1 U532 ( .A(KEYINPUT5), .B(KEYINPUT100), .Z(n440) );
  XNOR2_X1 U533 ( .A(G101), .B(G137), .ZN(n439) );
  XNOR2_X1 U534 ( .A(n443), .B(n442), .ZN(n660) );
  NAND2_X1 U535 ( .A1(n660), .A2(n465), .ZN(n444) );
  INV_X1 U536 ( .A(G472), .ZN(n658) );
  XNOR2_X2 U537 ( .A(n444), .B(n658), .ZN(n507) );
  INV_X1 U538 ( .A(KEYINPUT6), .ZN(n445) );
  INV_X1 U539 ( .A(n597), .ZN(n446) );
  NAND2_X1 U540 ( .A1(n506), .A2(n446), .ZN(n448) );
  XOR2_X1 U541 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n447) );
  XNOR2_X1 U542 ( .A(KEYINPUT96), .B(KEYINPUT17), .ZN(n449) );
  XNOR2_X1 U543 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U544 ( .A(n452), .B(n451), .ZN(n458) );
  NAND2_X1 U545 ( .A1(n453), .A2(G224), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n454), .B(KEYINPUT18), .ZN(n456) );
  XNOR2_X1 U547 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n458), .B(n457), .ZN(n461) );
  XNOR2_X1 U549 ( .A(KEYINPUT16), .B(G122), .ZN(n459) );
  XNOR2_X1 U550 ( .A(n460), .B(n459), .ZN(n767) );
  XNOR2_X1 U551 ( .A(n461), .B(n767), .ZN(n463) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n650) );
  NAND2_X1 U553 ( .A1(n650), .A2(n638), .ZN(n466) );
  NAND2_X1 U554 ( .A1(n465), .A2(n464), .ZN(n467) );
  NAND2_X1 U555 ( .A1(n467), .A2(G214), .ZN(n734) );
  NAND2_X1 U556 ( .A1(n601), .A2(n734), .ZN(n469) );
  INV_X1 U557 ( .A(KEYINPUT19), .ZN(n468) );
  NAND2_X1 U558 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U559 ( .A(n470), .B(KEYINPUT14), .ZN(n748) );
  NAND2_X1 U560 ( .A1(n769), .A2(G952), .ZN(n472) );
  NAND2_X1 U561 ( .A1(n345), .A2(G902), .ZN(n471) );
  NAND2_X1 U562 ( .A1(n472), .A2(n471), .ZN(n473) );
  AND2_X1 U563 ( .A1(n748), .A2(n473), .ZN(n570) );
  NAND2_X1 U564 ( .A1(n345), .A2(G898), .ZN(n474) );
  NAND2_X1 U565 ( .A1(n570), .A2(n474), .ZN(n475) );
  INV_X1 U566 ( .A(n528), .ZN(n476) );
  INV_X1 U567 ( .A(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n480), .B(n479), .ZN(n490) );
  XOR2_X1 U569 ( .A(n482), .B(n481), .Z(n488) );
  NAND2_X1 U570 ( .A1(G214), .A2(n483), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U572 ( .A(n486), .B(KEYINPUT11), .Z(n487) );
  XNOR2_X1 U573 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U574 ( .A(n490), .B(n489), .ZN(n641) );
  NOR2_X1 U575 ( .A1(G902), .A2(n641), .ZN(n492) );
  XNOR2_X1 U576 ( .A(KEYINPUT13), .B(G475), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n492), .B(n491), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT9), .B(G122), .Z(n495) );
  XNOR2_X1 U579 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U580 ( .A(n493), .B(n496), .ZN(n502) );
  INV_X1 U581 ( .A(G217), .ZN(n497) );
  OR2_X1 U582 ( .A1(n498), .A2(n497), .ZN(n500) );
  XOR2_X1 U583 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U584 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U585 ( .A(n502), .B(n501), .ZN(n677) );
  XNOR2_X1 U586 ( .A(G478), .B(n401), .ZN(n513) );
  NAND2_X1 U587 ( .A1(n512), .A2(n513), .ZN(n612) );
  XOR2_X1 U588 ( .A(KEYINPUT35), .B(KEYINPUT87), .Z(n503) );
  XNOR2_X2 U589 ( .A(n504), .B(n503), .ZN(n560) );
  AND2_X1 U590 ( .A1(KEYINPUT44), .A2(KEYINPUT90), .ZN(n505) );
  NAND2_X1 U591 ( .A1(n775), .A2(n505), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT101), .B(KEYINPUT31), .Z(n510) );
  INV_X1 U593 ( .A(n506), .ZN(n508) );
  NAND2_X1 U594 ( .A1(n730), .A2(n528), .ZN(n509) );
  XOR2_X1 U595 ( .A(n510), .B(n509), .Z(n703) );
  INV_X1 U596 ( .A(n513), .ZN(n511) );
  AND2_X1 U597 ( .A1(n512), .A2(n511), .ZN(n698) );
  OR2_X1 U598 ( .A1(n512), .A2(n511), .ZN(n704) );
  INV_X1 U599 ( .A(n704), .ZN(n695) );
  NOR2_X1 U600 ( .A1(n698), .A2(n695), .ZN(n739) );
  NOR2_X1 U601 ( .A1(n703), .A2(n739), .ZN(n524) );
  NOR2_X1 U602 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U603 ( .A(KEYINPUT103), .B(n514), .ZN(n737) );
  NOR2_X1 U604 ( .A1(n737), .A2(n721), .ZN(n515) );
  XNOR2_X1 U605 ( .A(n515), .B(KEYINPUT104), .ZN(n516) );
  XNOR2_X1 U606 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n518) );
  INV_X1 U607 ( .A(KEYINPUT66), .ZN(n517) );
  XNOR2_X1 U608 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U609 ( .A(n521), .ZN(n722) );
  NOR2_X1 U610 ( .A1(n346), .A2(n722), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n597), .A2(n522), .ZN(n523) );
  NOR2_X1 U612 ( .A1(n548), .A2(n523), .ZN(n688) );
  NAND2_X1 U613 ( .A1(n525), .A2(n725), .ZN(n527) );
  INV_X1 U614 ( .A(KEYINPUT98), .ZN(n526) );
  XNOR2_X2 U615 ( .A(n527), .B(n526), .ZN(n568) );
  NAND2_X1 U616 ( .A1(n568), .A2(n528), .ZN(n529) );
  XNOR2_X1 U617 ( .A(n529), .B(KEYINPUT99), .ZN(n530) );
  AND2_X1 U618 ( .A1(n530), .A2(n507), .ZN(n532) );
  NAND2_X1 U619 ( .A1(n698), .A2(n532), .ZN(n690) );
  NAND2_X1 U620 ( .A1(n531), .A2(n690), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n532), .A2(n695), .ZN(n693) );
  INV_X1 U622 ( .A(n693), .ZN(n533) );
  NOR2_X1 U623 ( .A1(n534), .A2(n533), .ZN(n537) );
  INV_X1 U624 ( .A(KEYINPUT90), .ZN(n535) );
  NAND2_X1 U625 ( .A1(n560), .A2(n535), .ZN(n536) );
  AND2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U627 ( .A(KEYINPUT44), .ZN(n540) );
  OR2_X1 U628 ( .A1(KEYINPUT65), .A2(n540), .ZN(n552) );
  OR2_X1 U629 ( .A1(n548), .A2(n346), .ZN(n542) );
  INV_X1 U630 ( .A(KEYINPUT106), .ZN(n541) );
  XNOR2_X1 U631 ( .A(n542), .B(n541), .ZN(n544) );
  AND2_X1 U632 ( .A1(n507), .A2(n722), .ZN(n543) );
  NAND2_X1 U633 ( .A1(n544), .A2(n543), .ZN(n656) );
  NAND2_X1 U634 ( .A1(n346), .A2(n722), .ZN(n545) );
  XNOR2_X1 U635 ( .A(n545), .B(KEYINPUT105), .ZN(n546) );
  NAND2_X1 U636 ( .A1(n546), .A2(n597), .ZN(n547) );
  OR2_X1 U637 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U638 ( .A(KEYINPUT32), .ZN(n549) );
  INV_X1 U639 ( .A(n777), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n656), .A2(n551), .ZN(n556) );
  AND2_X1 U641 ( .A1(n552), .A2(n556), .ZN(n555) );
  INV_X1 U642 ( .A(KEYINPUT65), .ZN(n564) );
  AND2_X1 U643 ( .A1(KEYINPUT91), .A2(n564), .ZN(n553) );
  NAND2_X1 U644 ( .A1(n560), .A2(n553), .ZN(n554) );
  NAND2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n558) );
  INV_X1 U646 ( .A(n556), .ZN(n561) );
  NAND2_X1 U647 ( .A1(n561), .A2(n564), .ZN(n557) );
  INV_X1 U648 ( .A(KEYINPUT91), .ZN(n559) );
  AND2_X1 U649 ( .A1(n560), .A2(n559), .ZN(n563) );
  AND2_X1 U650 ( .A1(n561), .A2(n540), .ZN(n562) );
  AND2_X1 U651 ( .A1(n564), .A2(KEYINPUT90), .ZN(n565) );
  OR2_X1 U652 ( .A1(KEYINPUT44), .A2(n565), .ZN(n566) );
  INV_X1 U653 ( .A(KEYINPUT45), .ZN(n567) );
  NOR2_X1 U654 ( .A1(n758), .A2(KEYINPUT2), .ZN(n634) );
  XNOR2_X1 U655 ( .A(n568), .B(KEYINPUT108), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n345), .A2(G900), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n570), .A2(n569), .ZN(n572) );
  INV_X1 U658 ( .A(KEYINPUT82), .ZN(n571) );
  XNOR2_X1 U659 ( .A(n572), .B(n571), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n573), .A2(n587), .ZN(n575) );
  INV_X1 U661 ( .A(KEYINPUT76), .ZN(n574) );
  XNOR2_X1 U662 ( .A(n575), .B(n574), .ZN(n580) );
  INV_X1 U663 ( .A(n734), .ZN(n576) );
  OR2_X1 U664 ( .A1(n507), .A2(n576), .ZN(n578) );
  INV_X1 U665 ( .A(KEYINPUT30), .ZN(n577) );
  XNOR2_X1 U666 ( .A(n578), .B(n577), .ZN(n579) );
  AND2_X2 U667 ( .A1(n580), .A2(n579), .ZN(n614) );
  INV_X1 U668 ( .A(KEYINPUT39), .ZN(n581) );
  INV_X1 U669 ( .A(KEYINPUT40), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U671 ( .A1(n737), .A2(n738), .ZN(n585) );
  XNOR2_X1 U672 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U675 ( .A1(n521), .A2(n589), .ZN(n590) );
  XOR2_X1 U676 ( .A(KEYINPUT70), .B(n590), .Z(n598) );
  NOR2_X1 U677 ( .A1(n598), .A2(n507), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(n403), .ZN(n592) );
  NAND2_X1 U679 ( .A1(n592), .A2(n525), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n593) );
  INV_X1 U681 ( .A(KEYINPUT88), .ZN(n594) );
  XNOR2_X1 U682 ( .A(n594), .B(KEYINPUT46), .ZN(n595) );
  XNOR2_X1 U683 ( .A(n596), .B(n595), .ZN(n620) );
  NOR2_X1 U684 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n599), .A2(n734), .ZN(n600) );
  INV_X1 U686 ( .A(n698), .ZN(n701) );
  NOR2_X1 U687 ( .A1(n600), .A2(n701), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n623), .A2(n601), .ZN(n602) );
  XOR2_X1 U689 ( .A(KEYINPUT36), .B(n602), .Z(n603) );
  NAND2_X1 U690 ( .A1(n603), .A2(n346), .ZN(n707) );
  XNOR2_X1 U691 ( .A(n707), .B(KEYINPUT89), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U693 ( .A(n739), .ZN(n608) );
  NOR2_X1 U694 ( .A1(n611), .A2(KEYINPUT47), .ZN(n609) );
  OR2_X1 U695 ( .A1(n610), .A2(n609), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n611), .A2(KEYINPUT47), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n655) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT85), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U701 ( .A(KEYINPUT48), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n622), .B(n621), .ZN(n632) );
  INV_X1 U703 ( .A(n346), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT43), .B(n625), .ZN(n626) );
  INV_X1 U706 ( .A(KEYINPUT107), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n628), .B(n627), .ZN(n774) );
  INV_X1 U708 ( .A(n629), .ZN(n630) );
  AND2_X1 U709 ( .A1(n630), .A2(n695), .ZN(n657) );
  NOR2_X1 U710 ( .A1(n774), .A2(n657), .ZN(n631) );
  INV_X1 U711 ( .A(KEYINPUT86), .ZN(n633) );
  XNOR2_X2 U712 ( .A(n635), .B(n633), .ZN(n664) );
  NAND2_X1 U713 ( .A1(n634), .A2(n664), .ZN(n637) );
  INV_X1 U714 ( .A(n758), .ZN(n709) );
  INV_X1 U715 ( .A(n635), .ZN(n710) );
  NAND2_X1 U716 ( .A1(n709), .A2(n710), .ZN(n714) );
  NAND2_X1 U717 ( .A1(n714), .A2(KEYINPUT2), .ZN(n636) );
  INV_X1 U718 ( .A(n638), .ZN(n639) );
  XNOR2_X1 U719 ( .A(KEYINPUT121), .B(KEYINPUT92), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n641), .B(KEYINPUT59), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U724 ( .A(KEYINPUT83), .B(KEYINPUT55), .Z(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT54), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U729 ( .A(n655), .B(G143), .ZN(G45) );
  XNOR2_X1 U730 ( .A(n656), .B(G110), .ZN(G12) );
  XOR2_X1 U731 ( .A(G134), .B(n657), .Z(G36) );
  XOR2_X1 U732 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G57) );
  BUF_X1 U736 ( .A(n664), .Z(n665) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(n670) );
  XOR2_X1 U738 ( .A(n670), .B(KEYINPUT125), .Z(n668) );
  XNOR2_X1 U739 ( .A(n665), .B(n668), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(n769), .ZN(n675) );
  XOR2_X1 U741 ( .A(G227), .B(n670), .Z(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(G900), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n672), .B(KEYINPUT126), .ZN(n673) );
  NAND2_X1 U744 ( .A1(n673), .A2(n345), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(G72) );
  NAND2_X1 U746 ( .A1(n680), .A2(G478), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n679), .A2(n686), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n680), .A2(G469), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT120), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(G54) );
  XOR2_X1 U755 ( .A(G101), .B(n688), .Z(n689) );
  XNOR2_X1 U756 ( .A(KEYINPUT114), .B(n689), .ZN(G3) );
  XNOR2_X1 U757 ( .A(G104), .B(n690), .ZN(G6) );
  XOR2_X1 U758 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n692) );
  XNOR2_X1 U759 ( .A(G107), .B(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(n694) );
  XOR2_X1 U761 ( .A(n694), .B(n693), .Z(G9) );
  XOR2_X1 U762 ( .A(G128), .B(KEYINPUT29), .Z(n697) );
  NAND2_X1 U763 ( .A1(n699), .A2(n695), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n697), .B(n696), .ZN(G30) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U766 ( .A(n700), .B(G146), .ZN(G48) );
  NOR2_X1 U767 ( .A1(n701), .A2(n703), .ZN(n702) );
  XOR2_X1 U768 ( .A(G113), .B(n702), .Z(G15) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U770 ( .A(G116), .B(n705), .Z(G18) );
  XOR2_X1 U771 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n706) );
  XNOR2_X1 U772 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U773 ( .A(G125), .B(n708), .ZN(G27) );
  NAND2_X1 U774 ( .A1(n710), .A2(KEYINPUT2), .ZN(n711) );
  NAND2_X1 U775 ( .A1(n709), .A2(n711), .ZN(n713) );
  INV_X1 U776 ( .A(n665), .ZN(n712) );
  NOR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n756) );
  AND2_X1 U778 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n714), .A2(n715), .ZN(n754) );
  NOR2_X1 U780 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n716) );
  NOR2_X1 U781 ( .A1(n345), .A2(n716), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n733), .A2(n717), .ZN(n718) );
  XNOR2_X1 U783 ( .A(n718), .B(KEYINPUT119), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n752) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U786 ( .A(KEYINPUT49), .B(n723), .Z(n724) );
  NAND2_X1 U787 ( .A1(n507), .A2(n724), .ZN(n728) );
  NOR2_X1 U788 ( .A1(n346), .A2(n725), .ZN(n726) );
  XNOR2_X1 U789 ( .A(n726), .B(KEYINPUT50), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U792 ( .A(KEYINPUT51), .B(n731), .Z(n732) );
  NOR2_X1 U793 ( .A1(n733), .A2(n732), .ZN(n745) );
  NOR2_X1 U794 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U795 ( .A1(n737), .A2(n736), .ZN(n742) );
  NOR2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U797 ( .A(KEYINPUT117), .B(n740), .Z(n741) );
  NOR2_X1 U798 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U799 ( .A1(n717), .A2(n743), .ZN(n744) );
  NOR2_X1 U800 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U801 ( .A(n746), .B(KEYINPUT118), .ZN(n747) );
  XNOR2_X1 U802 ( .A(n747), .B(KEYINPUT52), .ZN(n750) );
  NAND2_X1 U803 ( .A1(n748), .A2(G952), .ZN(n749) );
  NOR2_X1 U804 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U807 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U808 ( .A(KEYINPUT53), .B(n757), .ZN(G75) );
  BUF_X1 U809 ( .A(n758), .Z(n759) );
  NOR2_X1 U810 ( .A1(n759), .A2(n345), .ZN(n765) );
  NAND2_X1 U811 ( .A1(G224), .A2(n345), .ZN(n760) );
  XNOR2_X1 U812 ( .A(n760), .B(KEYINPUT61), .ZN(n761) );
  XNOR2_X1 U813 ( .A(KEYINPUT122), .B(n761), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n762), .A2(G898), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(KEYINPUT123), .ZN(n764) );
  NOR2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n773) );
  XNOR2_X1 U817 ( .A(n766), .B(KEYINPUT124), .ZN(n768) );
  XOR2_X1 U818 ( .A(n768), .B(n767), .Z(n771) );
  NOR2_X1 U819 ( .A1(n769), .A2(G898), .ZN(n770) );
  NOR2_X1 U820 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U821 ( .A(n773), .B(n772), .Z(G69) );
  XOR2_X1 U822 ( .A(G140), .B(n774), .Z(G42) );
  XOR2_X1 U823 ( .A(G122), .B(n775), .Z(G24) );
  XOR2_X1 U824 ( .A(G137), .B(n776), .Z(G39) );
  XOR2_X1 U825 ( .A(n777), .B(G119), .Z(G21) );
endmodule

