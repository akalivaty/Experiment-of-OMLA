//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  OR2_X1    g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n452), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n472), .B1(new_n481), .B2(G2105), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n464), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n470), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n468), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n485), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n468), .B(G138), .C1(KEYINPUT71), .C2(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(KEYINPUT71), .B2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n470), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  AND3_X1   g075(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(G651), .B1(new_n507), .B2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n501), .A2(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n508), .B1(new_n509), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n506), .A2(G51), .A3(G543), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(new_n521), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT74), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n503), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(new_n538), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n507), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n514), .A2(G90), .A3(new_n520), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n534), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n503), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G651), .B1(new_n507), .B2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n514), .A2(G81), .A3(new_n520), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(new_n514), .A2(new_n520), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n533), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G74), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n533), .B1(new_n503), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(G49), .B2(new_n507), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n521), .ZN(G288));
  AOI22_X1  g142(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n533), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(new_n570), .B1(G48), .B2(new_n507), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT75), .B1(new_n568), .B2(new_n533), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n556), .A2(G86), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n507), .A2(G47), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n521), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n533), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n503), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n507), .B2(G54), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n514), .A2(G92), .A3(new_n520), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n514), .A2(new_n520), .A3(new_n591), .A4(G92), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n590), .B1(new_n589), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n583), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n583), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G286), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g175(.A(G299), .B(KEYINPUT78), .Z(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G297));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G280));
  XOR2_X1   g178(.A(KEYINPUT79), .B(G559), .Z(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(G860), .B2(new_n604), .ZN(G148));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n478), .A2(new_n462), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  INV_X1    g188(.A(G123), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n485), .B2(new_n614), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n468), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n470), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n623), .ZN(G156));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2430), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT82), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  OR2_X1    g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G14), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n635), .B2(new_n638), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n639), .A2(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1981), .B(G1986), .ZN(new_n655));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT83), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n658), .A2(new_n659), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(new_n661), .ZN(new_n667));
  MUX2_X1   g242(.A(new_n667), .B(new_n666), .S(new_n657), .Z(new_n668));
  AOI21_X1  g243(.A(new_n655), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n665), .A2(new_n668), .A3(new_n655), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n673), .B1(new_n670), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n675), .B2(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G11), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT30), .B(G28), .Z(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G29), .ZN(new_n684));
  INV_X1    g259(.A(new_n622), .ZN(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G1966), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(G21), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G286), .B2(G16), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n684), .B(new_n687), .C1(new_n688), .C2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n688), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT93), .Z(new_n694));
  INV_X1    g269(.A(G1961), .ZN(new_n695));
  NOR2_X1   g270(.A1(G171), .A2(new_n689), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G5), .B2(new_n689), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n692), .B(new_n694), .C1(new_n695), .C2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G4), .A2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT88), .Z(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n595), .B2(new_n689), .ZN(new_n703));
  INV_X1    g278(.A(G1348), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(KEYINPUT23), .B1(new_n689), .B2(G20), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n707));
  AOI211_X1 g282(.A(new_n706), .B(new_n707), .C1(G299), .C2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT95), .B(G1956), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT96), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G34), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(G29), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G2084), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n550), .B2(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G1341), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n711), .A2(new_n712), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n686), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  INV_X1    g299(.A(G128), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G116), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n488), .B2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n686), .A2(G33), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n468), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n470), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(new_n686), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n717), .A2(new_n716), .B1(new_n743), .B2(G2072), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(G2072), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G1341), .B2(new_n720), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n722), .A2(new_n734), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2090), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n686), .A2(G32), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  INV_X1    g330(.A(G129), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n485), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n462), .A2(G105), .ZN(new_n758));
  INV_X1    g333(.A(G141), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n470), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n686), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT92), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G164), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G27), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n697), .A2(new_n695), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n751), .A2(new_n765), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n700), .A2(new_n705), .A3(new_n747), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G23), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n775));
  XNOR2_X1  g350(.A(G288), .B(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(new_n776), .B2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT33), .B(G1976), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(G6), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G305), .B2(new_n689), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT32), .B(G1981), .Z(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n689), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n689), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G1971), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G1971), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g366(.A(G290), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G16), .B2(G24), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n686), .A2(G25), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n488), .A2(G131), .ZN(new_n799));
  INV_X1    g374(.A(G119), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n468), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n485), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n686), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT85), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n797), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n791), .A2(new_n796), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n790), .A2(new_n811), .A3(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n811), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT36), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n810), .B(new_n817), .C1(new_n814), .C2(new_n813), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n773), .B1(new_n816), .B2(new_n818), .ZN(G311));
  INV_X1    g394(.A(new_n818), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n813), .A2(new_n814), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n817), .B1(new_n821), .B2(new_n810), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n772), .B1(new_n820), .B2(new_n822), .ZN(G150));
  OAI211_X1 g398(.A(G55), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n503), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n825), .B1(new_n828), .B2(G651), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n514), .A2(G93), .A3(new_n520), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n596), .A2(G559), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(KEYINPUT98), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n829), .A2(new_n837), .A3(new_n830), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n550), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n549), .A2(new_n831), .A3(KEYINPUT98), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n835), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT99), .Z(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n834), .B1(new_n846), .B2(new_n848), .ZN(G145));
  OR2_X1    g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n851));
  INV_X1    g426(.A(G142), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n851), .B1(new_n470), .B2(new_n852), .C1(new_n853), .C2(new_n485), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT104), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n611), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n804), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G164), .B(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(new_n732), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n496), .A2(new_n498), .ZN(new_n862));
  INV_X1    g437(.A(new_n493), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT102), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  NAND2_X1  g441(.A1(G164), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n732), .ZN(new_n869));
  INV_X1    g444(.A(new_n761), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n861), .B2(new_n869), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n737), .B2(new_n741), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n742), .A2(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n873), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n858), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n875), .B(new_n877), .C1(new_n872), .C2(new_n873), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n883), .A3(new_n871), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n857), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n881), .A2(KEYINPUT105), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G160), .B(KEYINPUT101), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G162), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n685), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n858), .B(new_n891), .C1(new_n876), .C2(new_n880), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n881), .B(new_n889), .C1(new_n895), .C2(new_n885), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n885), .A2(new_n895), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT40), .A4(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n886), .A2(new_n893), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n900), .A2(new_n904), .ZN(G395));
  NAND2_X1  g480(.A1(new_n831), .A2(new_n599), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n776), .B(G305), .ZN(new_n907));
  NAND2_X1  g482(.A1(G290), .A2(G166), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n579), .A2(G303), .A3(new_n581), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n908), .A2(new_n910), .ZN(new_n913));
  INV_X1    g488(.A(G305), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n776), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n912), .A2(new_n916), .A3(new_n918), .A4(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n606), .B(new_n841), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n595), .A2(new_n925), .A3(G299), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n589), .A2(new_n592), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT10), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G299), .A2(new_n925), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n557), .A2(KEYINPUT107), .A3(new_n559), .A4(new_n561), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n930), .A2(new_n587), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT41), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT41), .B1(new_n926), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT108), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT108), .B1(new_n926), .B2(new_n933), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n924), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n923), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n922), .A3(new_n921), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n906), .B1(new_n945), .B2(new_n599), .ZN(G295));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n906), .C1(new_n945), .C2(new_n599), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n599), .B1(new_n942), .B2(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(new_n906), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT110), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(G331));
  NAND2_X1  g527(.A1(new_n926), .A2(new_n933), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT41), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n829), .A2(new_n837), .A3(new_n830), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n837), .B1(new_n829), .B2(new_n830), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(new_n549), .ZN(new_n959));
  INV_X1    g534(.A(new_n840), .ZN(new_n960));
  NAND2_X1  g535(.A1(G301), .A2(G286), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(G301), .A2(G286), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n959), .A2(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n963), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(new_n839), .A3(new_n840), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n955), .A2(new_n956), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n841), .B(KEYINPUT112), .C1(new_n962), .C2(new_n963), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n926), .A3(new_n933), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n955), .A2(new_n975), .A3(new_n967), .A4(new_n956), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n969), .A2(new_n917), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n899), .ZN(new_n978));
  INV_X1    g553(.A(new_n967), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n938), .B2(new_n939), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n971), .A2(new_n972), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n980), .A2(KEYINPUT114), .B1(new_n936), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n979), .B(new_n983), .C1(new_n938), .C2(new_n939), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n917), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT115), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n976), .A2(new_n974), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n975), .B1(new_n936), .B2(new_n967), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n917), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n969), .A2(KEYINPUT113), .A3(new_n974), .A4(new_n976), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n978), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(KEYINPUT43), .C1(new_n978), .C2(new_n985), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n987), .A2(KEYINPUT44), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n994), .B2(new_n995), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n978), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n859), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n472), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n478), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1009));
  OAI211_X1 g584(.A(G40), .B(new_n1008), .C1(new_n1009), .C2(new_n468), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n761), .B(G1996), .ZN(new_n1014));
  INV_X1    g589(.A(G2067), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n732), .B(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n804), .B(new_n806), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n864), .A2(new_n1006), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n1010), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G164), .A2(G1384), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(G160), .A3(G40), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n571), .A2(new_n1030), .A3(new_n572), .A4(new_n573), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT118), .B(KEYINPUT49), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1028), .B(new_n1032), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n776), .A2(G1976), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1020), .B(new_n1023), .C1(new_n1011), .C2(new_n1025), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n1026), .B2(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  XOR2_X1   g619(.A(new_n1044), .B(KEYINPUT55), .Z(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1010), .B1(new_n1021), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n1006), .A4(new_n867), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1050));
  NAND3_X1  g625(.A1(new_n864), .A2(new_n1006), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1011), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1045), .C1(new_n1049), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1028), .A2(new_n1039), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1038), .A2(new_n1043), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1045), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n864), .A2(new_n1061), .A3(new_n1006), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1050), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(G164), .B2(G1384), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1011), .A3(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G2090), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1049), .A2(new_n1066), .A3(KEYINPUT119), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n1049), .B2(new_n1066), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1059), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1046), .B1(G164), .B2(G1384), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1011), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n688), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1051), .A2(new_n1011), .A3(new_n1052), .A4(new_n717), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1023), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1072), .B1(new_n1078), .B2(G286), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G286), .A2(G8), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT122), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1078), .B2(KEYINPUT121), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1083), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(G8), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n1072), .A3(new_n1080), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(KEYINPUT62), .A3(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1047), .A2(new_n1048), .A3(new_n768), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1092), .A2(new_n1093), .B1(new_n695), .B2(new_n1053), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1047), .A2(new_n1073), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1996), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1047), .A2(new_n1048), .A3(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1026), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n1103), .B2(new_n550), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1105), .B(new_n549), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1053), .A2(new_n704), .B1(new_n1022), .B2(new_n1015), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1053), .A2(new_n704), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1022), .A2(new_n1015), .ZN(new_n1111));
  AND4_X1   g686(.A1(KEYINPUT60), .A2(new_n1110), .A3(new_n595), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n595), .B1(new_n1108), .B2(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1047), .A2(new_n1048), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(G299), .B(KEYINPUT57), .Z(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1065), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1117), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1107), .A2(new_n1114), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n595), .B2(new_n1108), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G301), .B(KEYINPUT54), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n481), .A2(G2105), .B1(KEYINPUT123), .B2(new_n472), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1095), .A2(G40), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(KEYINPUT123), .C2(new_n472), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n859), .A2(new_n1006), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n1046), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1141), .B2(new_n1048), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1135), .A2(new_n1136), .B1(new_n1142), .B2(new_n1094), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1143), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1134), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1071), .B1(new_n1098), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G288), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1038), .A2(new_n1056), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1031), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1038), .A2(new_n1058), .A3(new_n1043), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1055), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1149), .A2(new_n1028), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1086), .A2(G286), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n1070), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(KEYINPUT63), .ZN(new_n1155));
  OAI21_X1  g730(.A(G8), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1155), .B(new_n1059), .C1(new_n1060), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1152), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1019), .B1(new_n1146), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1012), .A2(new_n795), .A3(new_n792), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT48), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1018), .A2(new_n1012), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n799), .A2(new_n803), .A3(new_n806), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1014), .A2(new_n1016), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n860), .A2(new_n1015), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1161), .A2(new_n1164), .B1(new_n1012), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT47), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1012), .A2(new_n1099), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(KEYINPUT124), .A3(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1016), .B(new_n761), .C1(new_n1172), .C2(G1996), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1012), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1170), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1174), .B(KEYINPUT46), .C1(new_n1012), .C2(new_n1099), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1170), .B(new_n1179), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1169), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT126), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1169), .B(new_n1187), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1159), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g765(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n1193), .A2(new_n679), .A3(new_n680), .ZN(new_n1194));
  XNOR2_X1  g768(.A(new_n1194), .B(KEYINPUT127), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1195), .B1(new_n902), .B2(new_n903), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1192), .A2(new_n1196), .ZN(G308));
  OAI221_X1 g771(.A(new_n1195), .B1(new_n903), .B2(new_n902), .C1(new_n1002), .C2(new_n1003), .ZN(G225));
endmodule


