//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(new_n201), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G116), .A2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n225), .B1(new_n202), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G68), .B2(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT65), .B(G77), .Z(new_n230));
  OAI211_X1 g0030(.A(new_n224), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n214), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n213), .B(new_n217), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G68), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n210), .B1(new_n214), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G77), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n211), .B2(G68), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n202), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT11), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT68), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT68), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n256), .B1(new_n268), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT12), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n265), .A2(G13), .A3(G20), .A4(new_n266), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n273), .B2(new_n249), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n264), .B1(new_n249), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n210), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n265), .A2(new_n284), .A3(new_n266), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(G238), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n226), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G97), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n294), .A2(new_n295), .A3(G232), .A4(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT73), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n288), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n302), .A2(KEYINPUT74), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT74), .B1(new_n302), .B2(new_n303), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n291), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n291), .C1(new_n304), .C2(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(KEYINPUT75), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(new_n312), .A3(KEYINPUT13), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n311), .A3(G169), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(G169), .A3(new_n313), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n307), .A2(G179), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n276), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n310), .A2(G200), .A3(new_n313), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n306), .B2(KEYINPUT13), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n276), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT77), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT70), .B(G58), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n207), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n255), .A2(KEYINPUT78), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G33), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT79), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n293), .A2(KEYINPUT79), .A3(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n333), .B(new_n211), .C1(new_n337), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G68), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n339), .A3(new_n340), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n333), .B1(new_n345), .B2(new_n211), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n332), .C1(new_n343), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n333), .A2(G20), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT3), .B1(new_n334), .B2(new_n336), .ZN(new_n350));
  INV_X1    g0150(.A(new_n295), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT3), .B(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n333), .B1(new_n353), .B2(G20), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n249), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n201), .B1(new_n329), .B2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(G159), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n211), .B1(new_n357), .B2(new_n261), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n348), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n347), .A2(new_n256), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT8), .A2(G58), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n329), .B2(KEYINPUT8), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n272), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n269), .B2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n226), .B2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n369), .A2(new_n344), .A3(new_n339), .A4(new_n340), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n286), .B1(new_n372), .B2(new_n303), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n287), .A2(KEYINPUT81), .A3(G232), .A4(new_n288), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G200), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n323), .A3(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT17), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT82), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n372), .A2(new_n303), .ZN(new_n386));
  AND4_X1   g0186(.A1(new_n323), .A2(new_n386), .A3(new_n285), .A4(new_n378), .ZN(new_n387));
  AOI21_X1  g0187(.A(G200), .B1(new_n373), .B2(new_n378), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n385), .B1(new_n366), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n360), .A4(new_n365), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n384), .B1(new_n392), .B2(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT80), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n360), .A2(new_n395), .A3(new_n365), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n379), .A2(G169), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n379), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT18), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n394), .A2(new_n402), .A3(new_n396), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n269), .A2(G50), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n203), .A2(G20), .ZN(new_n406));
  INV_X1    g0206(.A(G150), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n261), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n257), .B2(new_n362), .ZN(new_n409));
  INV_X1    g0209(.A(new_n256), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n405), .B1(G50), .B2(new_n272), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT9), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n285), .B1(new_n289), .B2(new_n226), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n353), .A2(G222), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g0216(.A(new_n416), .B(KEYINPUT69), .Z(new_n417));
  NAND2_X1  g0217(.A1(new_n353), .A2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G223), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(new_n230), .B2(new_n353), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n414), .B1(new_n421), .B2(new_n288), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  OAI211_X1 g0223(.A(G190), .B(new_n414), .C1(new_n421), .C2(new_n288), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n412), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT10), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT10), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n412), .A2(new_n427), .A3(new_n423), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n422), .A2(G179), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n411), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G77), .ZN(new_n434));
  INV_X1    g0234(.A(new_n230), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n270), .A2(new_n434), .B1(new_n435), .B2(new_n272), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n435), .A2(G20), .B1(new_n438), .B2(new_n257), .ZN(new_n439));
  XOR2_X1   g0239(.A(KEYINPUT8), .B(G58), .Z(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n260), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n410), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n353), .A2(G232), .A3(new_n415), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  INV_X1    g0245(.A(G238), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n444), .B1(new_n445), .B2(new_n353), .C1(new_n418), .C2(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n447), .A2(new_n303), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n285), .B1(new_n289), .B2(new_n229), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n443), .B1(new_n451), .B2(new_n431), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G179), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(G200), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(G190), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n454), .A2(new_n455), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n429), .A2(new_n433), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT72), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT72), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n429), .A2(new_n462), .A3(new_n433), .A4(new_n459), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n404), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n328), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n327), .A2(KEYINPUT77), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n352), .A2(new_n354), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G107), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n261), .A2(new_n434), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n221), .A2(new_n445), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT6), .A2(G97), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n476), .A2(KEYINPUT83), .A3(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT83), .B1(new_n476), .B2(G107), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n471), .B1(new_n479), .B2(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n410), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n272), .A2(G97), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n265), .A2(G33), .A3(new_n266), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n272), .A2(new_n410), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n485), .B2(G97), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n468), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(G20), .ZN(new_n489));
  INV_X1    g0289(.A(new_n471), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n445), .B1(new_n352), .B2(new_n354), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n256), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT84), .A3(new_n486), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n229), .A2(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n344), .A2(new_n339), .A3(new_n340), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT4), .A2(G244), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n294), .A2(new_n295), .A3(new_n499), .A4(new_n415), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n353), .A2(new_n502), .A3(new_n415), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n353), .A2(G250), .A3(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n303), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n265), .A2(G45), .A3(new_n266), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT5), .B(G41), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n280), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n288), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n222), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n507), .A2(new_n323), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(G200), .B1(new_n507), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n488), .B(new_n494), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n507), .A2(G179), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n496), .A2(new_n497), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n505), .A2(new_n504), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n503), .A4(new_n501), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n522), .B2(new_n303), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n431), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n493), .A2(new_n486), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n294), .A2(new_n295), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n211), .A2(G87), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n445), .A2(G20), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n334), .A2(new_n336), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n211), .A3(G116), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n339), .A2(new_n340), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n527), .A2(new_n219), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n537), .A2(new_n211), .A3(new_n344), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n536), .B2(new_n539), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n256), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n272), .A2(G107), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(G107), .B2(new_n485), .ZN(new_n548));
  XOR2_X1   g0348(.A(KEYINPUT91), .B(G294), .Z(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n534), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n222), .A2(G1698), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G250), .B2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n345), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n303), .B1(new_n509), .B2(new_n510), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n303), .B1(new_n554), .B2(G264), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n555), .A2(new_n323), .A3(new_n511), .ZN(new_n556));
  AOI21_X1  g0356(.A(G200), .B1(new_n555), .B2(new_n511), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n544), .B(new_n548), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n518), .A2(new_n526), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n504), .B(new_n211), .C1(G33), .C2(new_n221), .ZN(new_n560));
  INV_X1    g0360(.A(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n256), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n273), .A2(new_n561), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n272), .A2(new_n410), .A3(G116), .A4(new_n483), .ZN(new_n566));
  XOR2_X1   g0366(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(new_n256), .A3(new_n560), .A4(new_n562), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  MUX2_X1   g0369(.A(G257), .B(G264), .S(G1698), .Z(new_n570));
  NAND3_X1  g0370(.A1(new_n537), .A2(new_n344), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n528), .A2(G303), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n288), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G270), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n511), .B1(new_n513), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(KEYINPUT21), .B(G169), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n573), .A2(new_n575), .A3(new_n398), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n573), .A2(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  INV_X1    g0381(.A(new_n569), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n380), .C2(new_n580), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n569), .B(G169), .C1(new_n573), .C2(new_n575), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n579), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n555), .A2(new_n511), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n431), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n555), .A2(new_n398), .A3(new_n511), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n536), .A2(new_n539), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n540), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n410), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n548), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n591), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n537), .A2(new_n211), .A3(G68), .A4(new_n344), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n257), .A2(new_n600), .A3(G97), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n474), .A2(new_n219), .B1(new_n298), .B2(new_n211), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n410), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n438), .A2(new_n272), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n485), .A2(new_n438), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n534), .A2(G116), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n229), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G238), .B2(G1698), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n345), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n303), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n509), .A2(new_n280), .A3(KEYINPUT86), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n288), .A2(G274), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n508), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n303), .A2(new_n220), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n614), .A2(new_n617), .B1(new_n508), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n431), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n613), .A2(new_n619), .A3(new_n398), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(new_n619), .A3(G190), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(G200), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n484), .A2(new_n219), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n604), .A2(new_n605), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n613), .A2(new_n619), .A3(new_n629), .A4(G190), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n625), .A2(new_n626), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n598), .A2(new_n623), .A3(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n467), .A2(new_n559), .A3(new_n589), .A4(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n433), .ZN(new_n634));
  INV_X1    g0434(.A(new_n321), .ZN(new_n635));
  INV_X1    g0435(.A(new_n326), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n453), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n393), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n399), .A2(new_n366), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n634), .B1(new_n642), .B2(new_n429), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n608), .A2(new_n621), .A3(new_n622), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n631), .A2(new_n524), .A3(new_n623), .A4(new_n525), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT95), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n507), .A2(new_n515), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G169), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n488), .A2(new_n494), .B1(new_n649), .B2(new_n519), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n628), .A2(KEYINPUT92), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  NOR4_X1   g0453(.A1(new_n604), .A2(new_n627), .A3(new_n653), .A4(new_n605), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n626), .B(new_n624), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n650), .A2(new_n651), .A3(new_n655), .A4(new_n623), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n646), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n646), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n481), .A2(new_n468), .A3(new_n487), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT84), .B1(new_n493), .B2(new_n486), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n648), .A2(new_n380), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(G190), .B2(new_n648), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n662), .A2(new_n664), .B1(new_n525), .B2(new_n524), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT93), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n628), .B(KEYINPUT92), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n626), .A2(new_n624), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n644), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n665), .A2(new_n666), .A3(new_n669), .A4(new_n558), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n655), .A2(new_n623), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT93), .B1(new_n559), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n579), .B1(new_n587), .B2(new_n588), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT94), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n598), .ZN(new_n676));
  INV_X1    g0476(.A(new_n598), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT94), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n670), .A2(new_n672), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n659), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n643), .B1(new_n467), .B2(new_n680), .ZN(G369));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n211), .A2(G13), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n268), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G343), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n674), .B(new_n583), .C1(new_n582), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n673), .A2(new_n569), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT96), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n682), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n690), .B1(new_n596), .B2(new_n597), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n677), .B1(new_n558), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n598), .A2(new_n690), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n673), .A2(new_n688), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n698), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n215), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n474), .A2(new_n219), .A3(new_n561), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n281), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n209), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g0510(.A1(new_n646), .A2(new_n656), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT95), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n646), .A2(new_n647), .A3(new_n656), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n670), .A2(new_n672), .A3(new_n676), .A4(new_n678), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n690), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n623), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n651), .B1(new_n669), .B2(new_n650), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n671), .B(new_n559), .C1(new_n674), .C2(new_n598), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT29), .B(new_n688), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  OR4_X1    g0523(.A1(new_n559), .A2(new_n632), .A3(new_n589), .A4(new_n690), .ZN(new_n724));
  INV_X1    g0524(.A(new_n620), .ZN(new_n725));
  AND4_X1   g0525(.A1(new_n523), .A2(new_n725), .A3(new_n578), .A4(new_n555), .ZN(new_n726));
  OR2_X1    g0526(.A1(KEYINPUT97), .A2(KEYINPUT30), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n725), .A2(new_n580), .A3(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n648), .A3(new_n590), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n724), .A2(KEYINPUT31), .B1(new_n690), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT98), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n732), .A2(new_n736), .A3(KEYINPUT31), .A4(new_n690), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(G330), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n723), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n710), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n210), .B1(G20), .B2(new_n431), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n253), .A2(new_n283), .ZN(new_n748));
  INV_X1    g0548(.A(new_n345), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n705), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n283), .B2(new_n209), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n752), .B2(KEYINPUT99), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(KEYINPUT99), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n705), .A2(new_n528), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n755), .A2(G355), .B1(new_n561), .B2(new_n705), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n747), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n281), .B1(new_n683), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n706), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT100), .Z(new_n763));
  NOR2_X1   g0563(.A1(new_n323), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n323), .A2(new_n380), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G322), .A2(new_n766), .B1(new_n769), .B2(G326), .ZN(new_n770));
  INV_X1    g0570(.A(G329), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n323), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT101), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(G179), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n770), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n211), .A2(new_n323), .A3(new_n380), .A4(G179), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n528), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n774), .A2(G179), .A3(new_n380), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n764), .A2(new_n398), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n781), .B(new_n785), .C1(new_n549), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n763), .A2(new_n323), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n380), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n777), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT103), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT103), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT102), .B(G159), .Z(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n775), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT32), .Z(new_n802));
  AOI22_X1  g0602(.A1(G68), .A2(new_n794), .B1(new_n791), .B2(new_n435), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n783), .A2(new_n445), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n787), .A2(G97), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n805), .B(new_n353), .C1(new_n219), .C2(new_n779), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G50), .A2(new_n769), .B1(new_n766), .B2(new_n329), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n802), .A2(new_n803), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n797), .A2(new_n798), .A3(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n757), .B(new_n761), .C1(new_n810), .C2(new_n745), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n693), .A2(new_n694), .A3(new_n744), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n695), .A2(new_n760), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n693), .A2(new_n682), .A3(new_n694), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  AOI22_X1  g0618(.A1(G137), .A2(new_n769), .B1(new_n766), .B2(G143), .ZN(new_n819));
  INV_X1    g0619(.A(new_n794), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n820), .B2(new_n407), .C1(new_n792), .C2(new_n799), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  INV_X1    g0622(.A(new_n329), .ZN(new_n823));
  INV_X1    g0623(.A(new_n787), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n749), .B1(new_n779), .B2(new_n202), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n783), .A2(new_n249), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n776), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n822), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n353), .B1(new_n778), .B2(G107), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(new_n805), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n780), .B2(new_n768), .C1(new_n820), .C2(new_n784), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n783), .A2(new_n219), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n776), .A2(new_n789), .B1(new_n835), .B2(new_n765), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n792), .A2(new_n561), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n833), .A2(new_n834), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n745), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n745), .A2(new_n742), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n761), .B1(new_n434), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n458), .B1(new_n443), .B2(new_n688), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n453), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n453), .A2(new_n690), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n839), .B(new_n841), .C1(new_n846), .C2(new_n743), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n716), .A2(new_n846), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n688), .B(new_n846), .C1(new_n659), .C2(new_n679), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n739), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n761), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n848), .A2(new_n850), .A3(new_n739), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(G384));
  OR2_X1    g0654(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n212), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  NAND3_X1  g0658(.A1(new_n435), .A2(new_n209), .A3(new_n330), .ZN(new_n859));
  AOI211_X1 g0659(.A(G13), .B(new_n268), .C1(new_n859), .C2(new_n248), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n276), .A2(new_n690), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n321), .A2(new_n326), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n864));
  INV_X1    g0664(.A(new_n318), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n316), .B2(KEYINPUT14), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n315), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n276), .B(new_n690), .C1(new_n867), .C2(new_n636), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n732), .A2(new_n690), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n559), .A2(new_n632), .A3(new_n589), .A4(new_n690), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT31), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n845), .B1(new_n873), .B2(new_n734), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT108), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n394), .A2(new_n396), .A3(new_n687), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n640), .B1(new_n393), .B2(KEYINPUT106), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT17), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n390), .B2(new_n391), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n883), .B2(new_n384), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n879), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n879), .B(new_n639), .C1(new_n366), .C2(new_n389), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n879), .A2(new_n888), .A3(new_n390), .A4(new_n391), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n400), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n394), .A2(new_n891), .A3(new_n396), .A4(new_n399), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n878), .B1(new_n885), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n332), .B1(new_n343), .B2(new_n346), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n348), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n347), .A2(new_n256), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n365), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n687), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n404), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n399), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n392), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n893), .B2(new_n889), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(KEYINPUT38), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n877), .B1(new_n896), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n869), .A2(new_n910), .A3(new_n874), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n876), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n903), .A2(KEYINPUT38), .A3(new_n907), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n903), .B2(new_n907), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n869), .B(new_n874), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n873), .A2(new_n734), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n465), .A2(new_n466), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n392), .A2(KEYINPUT17), .ZN(new_n925));
  INV_X1    g0725(.A(new_n384), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(KEYINPUT106), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n641), .A3(new_n884), .ZN(new_n928));
  INV_X1    g0728(.A(new_n879), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n894), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n924), .B1(new_n931), .B2(new_n913), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n321), .A2(new_n690), .ZN(new_n933));
  INV_X1    g0733(.A(new_n914), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n641), .A2(new_n687), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n908), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n849), .A2(new_n844), .B1(new_n863), .B2(new_n868), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n849), .A2(new_n844), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n942), .A2(KEYINPUT104), .A3(new_n869), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n936), .B(new_n938), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n465), .A2(new_n717), .A3(new_n466), .A4(new_n722), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n643), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n923), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n268), .B2(new_n683), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n923), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n861), .B1(new_n949), .B2(new_n950), .ZN(G367));
  AOI22_X1  g0751(.A1(G143), .A2(new_n769), .B1(new_n775), .B2(G137), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n407), .B2(new_n765), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n353), .B1(new_n779), .B2(new_n823), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G68), .B2(new_n787), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n202), .B2(new_n792), .C1(new_n230), .C2(new_n783), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n953), .B(new_n956), .C1(new_n794), .C2(new_n800), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT113), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n780), .A2(new_n765), .B1(new_n768), .B2(new_n789), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n783), .A2(new_n221), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G317), .C2(new_n775), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n779), .B2(new_n561), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n787), .A2(G107), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n963), .A2(new_n345), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n794), .B2(new_n549), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n961), .B(new_n967), .C1(new_n784), .C2(new_n792), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n958), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n745), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n750), .A2(new_n238), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n747), .B1(new_n705), .B2(new_n438), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n761), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n744), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n667), .A2(new_n688), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n669), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n623), .B2(new_n976), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n971), .B(new_n974), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n665), .B1(new_n662), .B2(new_n688), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n650), .A2(new_n690), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n702), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n677), .B1(new_n525), .B2(new_n524), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n986), .C1(new_n987), .C2(new_n690), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT109), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n978), .B(KEYINPUT43), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n989), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n695), .A2(new_n699), .A3(new_n983), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n740), .ZN(new_n997));
  INV_X1    g0797(.A(new_n703), .ZN(new_n998));
  INV_X1    g0798(.A(new_n983), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT110), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT110), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n703), .A2(new_n1001), .A3(new_n983), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n999), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n703), .B2(new_n983), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n700), .A2(KEYINPUT112), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n700), .A2(KEYINPUT112), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT45), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1014));
  OAI211_X1 g0814(.A(KEYINPUT112), .B(new_n700), .C1(new_n1014), .C2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n699), .B(new_n701), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n695), .B2(KEYINPUT111), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n695), .B(KEYINPUT111), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n1017), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n997), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n706), .B(KEYINPUT41), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n758), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n980), .B1(new_n996), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(G387));
  NAND2_X1  g0825(.A1(new_n1020), .A2(new_n740), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n706), .B(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT116), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(KEYINPUT116), .A3(new_n1027), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n740), .C2(new_n1020), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n755), .A2(new_n707), .B1(new_n445), .B2(new_n705), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n243), .A2(new_n283), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n440), .A2(new_n202), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n707), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n283), .C1(new_n249), .C2(new_n434), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n750), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1033), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n761), .B1(new_n1040), .B2(new_n746), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n699), .B2(new_n975), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n202), .A2(new_n765), .B1(new_n768), .B2(new_n357), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1043), .B(new_n960), .C1(G150), .C2(new_n775), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n824), .A2(new_n437), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n749), .B1(new_n230), .B2(new_n779), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G68), .C2(new_n791), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1047), .C1(new_n363), .C2(new_n820), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n749), .B1(new_n775), .B2(G326), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n766), .B1(new_n769), .B2(G322), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n820), .B2(new_n789), .C1(new_n780), .C2(new_n792), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n787), .A2(G283), .B1(new_n778), .B2(new_n549), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT49), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1049), .B1(new_n561), .B2(new_n783), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1048), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1042), .B1(new_n1060), .B2(new_n745), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT114), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1020), .B2(new_n759), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1032), .A2(new_n1063), .ZN(G393));
  NAND3_X1  g0864(.A1(new_n1016), .A2(new_n740), .A3(new_n1020), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1026), .A2(new_n1015), .A3(new_n1013), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n1027), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n999), .A2(new_n744), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n746), .B1(new_n221), .B2(new_n215), .C1(new_n751), .C2(new_n247), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n760), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n766), .B1(new_n769), .B2(G317), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  OAI221_X1 g0872(.A(new_n528), .B1(new_n779), .B2(new_n784), .C1(new_n824), .C2(new_n561), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1073), .B(new_n804), .C1(G322), .C2(new_n775), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G294), .A2(new_n791), .B1(new_n794), .B2(G303), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n824), .A2(new_n434), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n791), .B2(new_n440), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n202), .B2(new_n820), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT117), .Z(new_n1080));
  AOI211_X1 g0880(.A(new_n345), .B(new_n834), .C1(G68), .C2(new_n778), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n407), .A2(new_n768), .B1(new_n765), .B2(new_n357), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n775), .A2(G143), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1070), .B1(new_n1086), .B2(new_n745), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1016), .A2(new_n759), .B1(new_n1068), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1067), .A2(new_n1088), .ZN(G390));
  INV_X1    g0889(.A(new_n840), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n760), .B1(new_n362), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n528), .B1(new_n779), .B2(new_n219), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n826), .A2(new_n1077), .A3(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n221), .B2(new_n792), .C1(new_n445), .C2(new_n820), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G116), .A2(new_n766), .B1(new_n769), .B2(G283), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n835), .B2(new_n776), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G128), .A2(new_n769), .B1(new_n775), .B2(G125), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n202), .B2(new_n783), .C1(new_n828), .C2(new_n765), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n778), .A2(G150), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT53), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n794), .A2(G137), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n791), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n528), .B1(new_n787), .B2(G159), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1101), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1094), .A2(new_n1096), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n745), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n932), .A2(new_n935), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n743), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n942), .A2(new_n869), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n321), .B2(new_n690), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1109), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n863), .A2(new_n868), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n688), .B1(new_n720), .B2(new_n721), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n843), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n844), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n869), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n933), .B1(new_n896), .B2(new_n908), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(G330), .B(new_n846), .C1(new_n733), .C2(new_n738), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n869), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1114), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1113), .A2(new_n1109), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n874), .A2(G330), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1115), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1126), .A2(new_n869), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n942), .B1(new_n1134), .B2(new_n1131), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1130), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1119), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1127), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n682), .B1(new_n873), .B2(new_n734), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n465), .A2(new_n466), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n945), .A2(new_n643), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT119), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT119), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n945), .A2(new_n1142), .A3(new_n643), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1027), .B1(new_n1133), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1133), .A2(new_n1147), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1111), .B1(new_n758), .B2(new_n1133), .C1(new_n1148), .C2(new_n1149), .ZN(G378));
  OAI21_X1  g0950(.A(new_n760), .B1(G50), .B2(new_n1090), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n791), .A2(new_n438), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n775), .A2(G283), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n435), .A2(new_n778), .B1(new_n787), .B2(G68), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G107), .A2(new_n766), .B1(new_n769), .B2(G116), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n749), .A2(G41), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n823), .C2(new_n783), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(G97), .C2(new_n794), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT58), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G132), .A2(new_n794), .B1(new_n791), .B2(G137), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1103), .A2(new_n778), .B1(G150), .B2(new_n787), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G125), .A2(new_n769), .B1(new_n766), .B2(G128), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n255), .B(new_n282), .C1(new_n783), .C2(new_n799), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G124), .B2(new_n775), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1159), .A2(KEYINPUT58), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1157), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1160), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1151), .B1(new_n1173), .B2(new_n745), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n429), .A2(new_n433), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n411), .A2(new_n687), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1174), .B1(new_n1179), .B2(new_n743), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT121), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n682), .B1(new_n915), .B2(new_n916), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n912), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1179), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n912), .A2(new_n1183), .A3(new_n1179), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n943), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n913), .A2(new_n914), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT104), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1112), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n937), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1186), .A2(new_n1187), .B1(new_n1192), .B2(new_n936), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n912), .A2(new_n1183), .A3(new_n1179), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1179), .B1(new_n912), .B2(new_n1183), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n944), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1182), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1186), .A2(new_n936), .A3(new_n1192), .A4(new_n1187), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n944), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1181), .B1(new_n1201), .B2(new_n759), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1140), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1133), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1027), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1207), .B2(new_n1210), .ZN(G375));
  XNOR2_X1  g1011(.A(new_n1022), .B(KEYINPUT122), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1204), .B2(new_n1140), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(new_n1203), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n743), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT123), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n760), .B1(G68), .B2(new_n1090), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n783), .A2(new_n434), .B1(new_n784), .B2(new_n765), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G294), .B2(new_n769), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n791), .A2(G107), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n794), .A2(G116), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n528), .B1(new_n779), .B2(new_n221), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1045), .B(new_n1223), .C1(G303), .C2(new_n775), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n749), .B1(new_n779), .B2(new_n357), .C1(new_n202), .C2(new_n824), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n775), .A2(G128), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n783), .B2(new_n823), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G150), .C2(new_n791), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT124), .Z(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n769), .B1(new_n766), .B2(G137), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n794), .A2(new_n1103), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1218), .B1(new_n1234), .B2(new_n745), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1217), .A2(new_n1235), .B1(new_n1140), .B2(new_n759), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1215), .A2(new_n1236), .ZN(G381));
  OR2_X1    g1037(.A1(G390), .A2(G384), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1032), .A2(new_n817), .A3(new_n1063), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(G387), .A2(new_n1238), .A3(G381), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G375), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1111), .B1(new_n1133), .B2(new_n758), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G343), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G213), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1241), .A2(new_n1244), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(new_n1249), .A3(G213), .ZN(G409));
  OAI211_X1 g1050(.A(G378), .B(new_n1202), .C1(new_n1207), .C2(new_n1210), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1181), .B1(new_n1208), .B2(new_n759), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT121), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT121), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1206), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1252), .B1(new_n1255), .B2(new_n1212), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1244), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1247), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1248), .A2(G2897), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT126), .Z(new_n1261));
  NOR2_X1   g1061(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1140), .B1(new_n1146), .B2(new_n1144), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT60), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1027), .B(new_n1147), .C1(new_n1264), .C2(KEYINPUT60), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1236), .B(new_n1263), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n1262), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1214), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1273), .A2(new_n1265), .A3(new_n1027), .A4(new_n1147), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1274), .B2(new_n1236), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1261), .B1(new_n1269), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1261), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1274), .A2(new_n1236), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1268), .B(new_n1277), .C1(new_n1278), .C2(new_n1271), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1259), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1239), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n817), .B1(new_n1032), .B2(new_n1063), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1024), .B2(G390), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1024), .A2(G390), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1024), .A2(G390), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1288), .A2(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1024), .A2(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1239), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1024), .A2(G390), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1248), .B1(new_n1251), .B2(new_n1257), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1281), .A2(new_n1285), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1299), .A2(new_n1302), .A3(new_n1283), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1299), .B2(new_n1283), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1301), .B1(new_n1308), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1109(.A1(new_n1298), .A2(new_n1283), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1292), .A2(new_n1297), .A3(new_n1284), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G375), .B(G378), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1312), .B(new_n1313), .ZN(G402));
endmodule


