//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G217), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G122), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(G116), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(G107), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT68), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT68), .A2(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(G143), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT93), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(KEYINPUT93), .B(G143), .C1(new_n198), .C2(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n207), .A2(KEYINPUT13), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT93), .B1(new_n212), .B2(G143), .ZN(new_n213));
  INV_X1    g027(.A(new_n203), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT94), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n204), .A2(KEYINPUT94), .A3(new_n211), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(KEYINPUT13), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI211_X1 g034(.A(new_n197), .B(new_n210), .C1(new_n220), .C2(G134), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT14), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n195), .B1(new_n193), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT95), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n194), .A2(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g039(.A(G107), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n196), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n205), .B1(new_n204), .B2(new_n208), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(new_n228), .C1(new_n210), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n191), .B1(new_n221), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(G134), .ZN(new_n233));
  INV_X1    g047(.A(new_n197), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n209), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n230), .A3(new_n190), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(KEYINPUT96), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT96), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n239), .A3(new_n230), .A4(new_n190), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT15), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G478), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(G478), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n237), .A2(new_n238), .A3(new_n240), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G475), .ZN(new_n248));
  XNOR2_X1  g062(.A(G113), .B(G122), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n249), .A2(G104), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(G104), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G214), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G131), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n253), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G125), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT89), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT19), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT16), .ZN(new_n273));
  INV_X1    g087(.A(G140), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(G125), .ZN(new_n276));
  INV_X1    g090(.A(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G140), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n279), .B2(new_n273), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(new_n271), .ZN(new_n281));
  INV_X1    g095(.A(new_n261), .ZN(new_n282));
  AOI21_X1  g096(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n283));
  OAI21_X1  g097(.A(G131), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT88), .A3(new_n262), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n265), .A2(new_n272), .A3(new_n281), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT18), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n258), .B(new_n261), .C1(new_n287), .C2(new_n259), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n279), .A2(G146), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n266), .A2(new_n271), .ZN(new_n290));
  OAI221_X1 g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .C1(new_n284), .C2(new_n287), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n252), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n293), .A3(new_n262), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n271), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n294), .A2(new_n281), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT90), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n250), .A2(new_n298), .A3(new_n251), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n250), .B2(new_n251), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n297), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n248), .B(new_n238), .C1(new_n292), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT91), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(KEYINPUT20), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n292), .A2(new_n302), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n248), .A4(new_n238), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT20), .A3(new_n304), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n252), .B1(new_n297), .B2(new_n291), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n238), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(G475), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n247), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n255), .A2(G952), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(G234), .B2(G237), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  NAND2_X1  g136(.A1(G234), .A2(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G902), .A3(G953), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G472), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n260), .A2(G210), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT27), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT26), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(KEYINPUT2), .A2(G113), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT2), .A2(G113), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G116), .ZN(new_n339));
  INV_X1    g153(.A(G116), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G119), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n339), .B2(new_n341), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n335), .A2(new_n339), .A3(new_n341), .A4(new_n336), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT71), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n337), .C1(new_n343), .C2(new_n344), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT67), .ZN(new_n353));
  XNOR2_X1  g167(.A(G134), .B(G137), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n259), .ZN(new_n355));
  INV_X1    g169(.A(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G134), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n205), .A2(G137), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT67), .A3(G131), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(KEYINPUT11), .A3(G134), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(new_n358), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT11), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT66), .B(new_n364), .C1(new_n205), .C2(G137), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT66), .B1(new_n357), .B2(new_n364), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n363), .B(new_n259), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT72), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(new_n361), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n271), .A2(G143), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n271), .A2(G143), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(KEYINPUT65), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n271), .A3(G143), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n374), .A2(new_n375), .A3(G128), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n257), .A2(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n375), .B1(G143), .B2(new_n271), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n212), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n370), .A2(new_n371), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G131), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n368), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT0), .A2(G128), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(KEYINPUT64), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT65), .B1(new_n257), .B2(G146), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n257), .A2(G146), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n377), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n390), .A2(KEYINPUT0), .A3(G128), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT0), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n380), .A2(new_n389), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(KEYINPUT64), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT30), .B1(new_n385), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n383), .A2(new_n368), .A3(new_n361), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n352), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n361), .A2(new_n368), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT72), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n383), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n352), .A3(new_n399), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n334), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(KEYINPUT28), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(new_n415), .A3(new_n352), .A4(new_n399), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n399), .A2(new_n402), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n351), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n333), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n413), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n334), .A2(new_n413), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n352), .B1(new_n409), .B2(new_n399), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n414), .B2(new_n416), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n328), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G472), .A2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n403), .B1(new_n409), .B2(new_n399), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n351), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n431), .A2(new_n410), .A3(new_n333), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT31), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n417), .A2(new_n419), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n334), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n410), .A3(new_n333), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT31), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n428), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n426), .B1(new_n438), .B2(KEYINPUT32), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n334), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n431), .A2(new_n433), .A3(new_n410), .A4(new_n333), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n437), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n427), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n281), .A2(new_n295), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT74), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT74), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT23), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n451), .B(new_n453), .C1(new_n338), .C2(G128), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT23), .B(G119), .C1(new_n198), .C2(new_n199), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n338), .A2(G128), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT75), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT75), .A4(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(G110), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n212), .A2(G119), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n456), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT24), .B(G110), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n449), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n289), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n457), .A2(G110), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n281), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(G221), .A2(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT76), .B1(new_n470), .B2(G953), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(new_n255), .A3(G221), .A4(G234), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT22), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n471), .B2(new_n473), .ZN(new_n477));
  OR3_X1    g291(.A1(new_n476), .A2(new_n356), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n356), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n465), .A2(new_n469), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n465), .B2(new_n469), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n481), .A2(new_n482), .A3(G902), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n448), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n189), .B1(G234), .B2(new_n238), .ZN(new_n486));
  INV_X1    g300(.A(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n465), .A2(new_n469), .A3(new_n480), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n238), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n486), .A2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(KEYINPUT78), .A3(new_n495), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n439), .A2(new_n447), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(G110), .B(G122), .Z(new_n503));
  INV_X1    g317(.A(G104), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT3), .B1(new_n504), .B2(G107), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT3), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n227), .A3(G104), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(G107), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n332), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n510), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n351), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n339), .A2(new_n341), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT69), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n338), .A3(G116), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(G113), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n515), .A2(new_n516), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n227), .A2(G104), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n504), .A2(G107), .ZN(new_n526));
  OAI21_X1  g340(.A(G101), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n509), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT82), .B1(new_n514), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n503), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n514), .A2(new_n530), .ZN(new_n534));
  INV_X1    g348(.A(new_n503), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n398), .A2(G125), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n383), .A2(new_n277), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT84), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G224), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n543), .B(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n533), .A2(new_n548), .A3(KEYINPUT6), .A4(new_n536), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n538), .A2(new_n546), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  OR3_X1    g364(.A1(new_n524), .A2(KEYINPUT85), .A3(new_n529), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n523), .B1(new_n521), .B2(new_n517), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n348), .A2(new_n529), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT85), .B1(new_n524), .B2(new_n529), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n503), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n545), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n534), .A2(new_n535), .B1(new_n541), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n541), .A2(new_n561), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(KEYINPUT86), .A3(new_n556), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n550), .A2(new_n238), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n567), .B(KEYINPUT87), .Z(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n550), .A2(new_n238), .A3(new_n567), .A4(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n502), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G469), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n573));
  OAI21_X1  g387(.A(G128), .B1(new_n381), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n372), .A2(new_n573), .A3(KEYINPUT1), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n393), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n528), .B1(new_n577), .B2(new_n378), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n378), .A2(new_n528), .A3(new_n382), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n388), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT12), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n388), .B(KEYINPUT12), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n509), .A2(new_n527), .A3(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n383), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n383), .A2(KEYINPUT80), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n578), .A2(KEYINPUT10), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n387), .A2(new_n368), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n513), .A2(new_n398), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(G110), .B(G140), .Z(new_n595));
  INV_X1    g409(.A(G227), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(G953), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n595), .B(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n584), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n589), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT80), .B1(new_n383), .B2(new_n585), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n398), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n510), .A2(G101), .A3(new_n511), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n509), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n603), .A2(new_n606), .B1(new_n578), .B2(KEYINPUT10), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n388), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n598), .B1(new_n608), .B2(new_n594), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n572), .B(new_n238), .C1(new_n599), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(G469), .A2(G902), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n594), .A3(new_n598), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n584), .A2(new_n594), .ZN(new_n613));
  OAI211_X1 g427(.A(G469), .B(new_n612), .C1(new_n613), .C2(new_n598), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT81), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n327), .A2(new_n500), .A3(new_n571), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NAND2_X1  g437(.A1(new_n498), .A2(new_n499), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n238), .B1(new_n442), .B2(new_n443), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n444), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n620), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n237), .A2(new_n633), .A3(new_n240), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n232), .A2(KEYINPUT33), .A3(new_n236), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n241), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n316), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n501), .B1(new_n570), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n567), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n566), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n570), .A2(new_n642), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n632), .A2(new_n326), .A3(new_n641), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND2_X1  g465(.A1(new_n246), .A2(new_n317), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT99), .B1(new_n652), .B2(new_n326), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n246), .A2(new_n654), .A3(new_n325), .A4(new_n317), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n648), .B(new_n632), .C1(new_n653), .C2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT35), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G107), .ZN(G9));
  INV_X1    g472(.A(new_n480), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT36), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n465), .A2(new_n469), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n494), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n491), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n318), .A2(new_n326), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n626), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n438), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n571), .A3(new_n621), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT37), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G110), .ZN(G12));
  AOI22_X1  g485(.A1(new_n439), .A2(new_n447), .B1(new_n618), .B2(new_n620), .ZN(new_n672));
  INV_X1    g486(.A(new_n643), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n645), .A2(new_n642), .A3(new_n570), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n324), .A2(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n321), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n246), .A2(new_n317), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n665), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n676), .B(KEYINPUT39), .Z(new_n681));
  OAI21_X1  g495(.A(KEYINPUT40), .B1(new_n630), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n334), .B1(new_n411), .B2(new_n423), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n436), .A2(new_n683), .A3(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(G472), .A2(G902), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n447), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(KEYINPUT32), .B(new_n427), .C1(new_n442), .C2(new_n443), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(KEYINPUT100), .B2(new_n686), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT101), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n686), .A2(KEYINPUT100), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n438), .B2(KEYINPUT32), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n444), .A2(new_n446), .B1(new_n686), .B2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n697));
  INV_X1    g511(.A(new_n681), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n621), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n682), .A2(new_n691), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n247), .A2(new_n317), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT38), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n569), .A2(new_n702), .A3(new_n570), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n569), .B2(new_n570), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n501), .B(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n700), .A2(new_n705), .A3(new_n664), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n257), .ZN(G45));
  NAND3_X1  g521(.A1(new_n640), .A2(new_n316), .A3(new_n676), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n665), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(new_n641), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n599), .A2(new_n609), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n238), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n610), .ZN(new_n716));
  INV_X1    g530(.A(new_n616), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n326), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n647), .A2(new_n500), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT41), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G113), .ZN(G15));
  NAND2_X1  g535(.A1(new_n653), .A2(new_n655), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n716), .A2(new_n717), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n647), .A2(new_n722), .A3(new_n500), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND2_X1  g539(.A1(new_n439), .A2(new_n447), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n647), .A2(new_n666), .A3(new_n726), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  OAI21_X1  g542(.A(new_n441), .B1(new_n333), .B2(new_n424), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n427), .B1(new_n443), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n667), .A2(new_n731), .A3(new_n496), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n647), .A2(new_n701), .A3(new_n718), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  AOI21_X1  g548(.A(G902), .B1(new_n435), .B2(new_n437), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n664), .B(new_n730), .C1(new_n735), .C2(new_n328), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n708), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n673), .A3(new_n674), .A4(new_n723), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  OR2_X1    g553(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n496), .B1(new_n740), .B2(new_n439), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n569), .A2(new_n501), .A3(new_n570), .ZN(new_n742));
  INV_X1    g556(.A(new_n617), .ZN(new_n743));
  INV_X1    g557(.A(new_n708), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n426), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n689), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n438), .A2(new_n445), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n624), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n569), .A2(new_n501), .A3(new_n570), .A4(new_n743), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n708), .A2(KEYINPUT42), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n745), .A2(KEYINPUT42), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NOR3_X1   g568(.A1(new_n749), .A2(new_n750), .A3(new_n677), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n205), .ZN(G36));
  NAND2_X1  g570(.A1(new_n640), .A2(new_n317), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n316), .B1(new_n638), .B2(new_n639), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g578(.A(new_n668), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT104), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n758), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n765), .A3(new_n664), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n569), .A2(new_n501), .A3(new_n570), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n612), .B1(new_n613), .B2(new_n598), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n612), .C1(new_n613), .C2(new_n598), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(G469), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n611), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n611), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n610), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n616), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n698), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n616), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT102), .B1(new_n785), .B2(new_n681), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n771), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n668), .B1(new_n763), .B2(KEYINPUT104), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n664), .A4(new_n767), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n770), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  AND2_X1   g605(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n726), .A2(new_n624), .A3(new_n708), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n742), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n679), .A2(new_n710), .A3(new_n738), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n673), .A2(new_n674), .A3(new_n701), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n665), .B(new_n676), .C1(new_n688), .C2(new_n690), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n799), .A2(new_n800), .A3(new_n617), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  INV_X1    g617(.A(new_n800), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n647), .A3(new_n743), .A4(new_n701), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n647), .B(new_n672), .C1(new_n678), .C2(new_n709), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n738), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n802), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n803), .B1(new_n802), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n641), .A2(new_n652), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n631), .A2(new_n325), .A3(new_n571), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n724), .A3(new_n733), .A4(new_n669), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n727), .A2(new_n719), .A3(new_n622), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n750), .A2(new_n708), .A3(new_n736), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n755), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT105), .ZN(new_n821));
  INV_X1    g635(.A(new_n676), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n246), .A2(new_n821), .A3(new_n316), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n771), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n318), .B2(new_n822), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n664), .A3(new_n825), .A4(new_n672), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT106), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n755), .ZN(new_n829));
  INV_X1    g643(.A(new_n819), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n826), .A3(new_n830), .A4(KEYINPUT106), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n818), .A2(new_n828), .A3(new_n753), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n811), .A2(new_n813), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n802), .A2(new_n808), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT107), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT107), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n802), .A2(new_n836), .A3(new_n808), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n753), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n839), .A2(new_n827), .A3(new_n816), .A4(new_n817), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n813), .B1(new_n811), .B2(new_n832), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  INV_X1    g662(.A(new_n763), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n771), .A2(new_n717), .A3(new_n716), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n320), .A4(new_n741), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n691), .A2(new_n696), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n850), .ZN(new_n854));
  INV_X1    g668(.A(new_n640), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n321), .B1(new_n498), .B2(new_n499), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n317), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n849), .A3(new_n320), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n736), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT112), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n320), .A2(new_n732), .A3(new_n758), .A4(new_n762), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n502), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n703), .A2(new_n704), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n723), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n865), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n502), .A4(new_n862), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n862), .A2(new_n742), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n715), .A2(new_n717), .A3(new_n610), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n792), .B2(new_n793), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n859), .B2(KEYINPUT112), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n647), .A2(new_n723), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n862), .A2(new_n877), .B1(new_n878), .B2(new_n319), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n854), .A2(new_n712), .A3(new_n856), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n880), .C1(new_n878), .C2(new_n319), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n870), .A2(new_n876), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n873), .B(KEYINPUT110), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n872), .B1(new_n794), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n871), .B1(new_n888), .B2(new_n859), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT111), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(KEYINPUT111), .B(new_n871), .C1(new_n888), .C2(new_n859), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n847), .A2(new_n848), .A3(new_n852), .A4(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n842), .A3(new_n852), .A4(new_n846), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT115), .ZN(new_n896));
  OR2_X1    g710(.A1(G952), .A2(G953), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n501), .A2(new_n853), .A3(new_n616), .A4(new_n760), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n716), .A2(KEYINPUT49), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n496), .B1(new_n716), .B2(KEYINPUT49), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n864), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n255), .A2(G952), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n538), .A2(new_n547), .A3(new_n549), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n546), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT116), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT55), .Z(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n238), .B1(new_n843), .B2(new_n845), .ZN(new_n910));
  AOI211_X1 g724(.A(KEYINPUT56), .B(new_n909), .C1(new_n910), .C2(new_n568), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n843), .A2(new_n845), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n916), .A3(G210), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n904), .B(new_n911), .C1(new_n918), .C2(new_n909), .ZN(G51));
  XOR2_X1   g733(.A(new_n611), .B(KEYINPUT57), .Z(new_n920));
  AND3_X1   g734(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n920), .C1(new_n921), .C2(new_n922), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n713), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n776), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n910), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n904), .B1(new_n927), .B2(new_n929), .ZN(G54));
  INV_X1    g744(.A(KEYINPUT58), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT119), .B1(new_n931), .B2(new_n248), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n931), .A2(new_n248), .A3(KEYINPUT119), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n910), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n306), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n904), .ZN(G60));
  NAND2_X1  g752(.A1(new_n634), .A2(new_n635), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n847), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n904), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n939), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n921), .B2(new_n922), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n843), .B2(new_n845), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(new_n493), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n950), .A2(new_n952), .A3(new_n662), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n950), .B2(new_n662), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n943), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n949), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n912), .A2(new_n662), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n950), .A2(new_n952), .A3(new_n662), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n943), .A4(new_n951), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n957), .A2(new_n963), .ZN(G66));
  INV_X1    g778(.A(new_n322), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n965), .B2(new_n544), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n818), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n905), .B1(G898), .B2(new_n255), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  NOR2_X1   g783(.A1(new_n429), .A2(new_n430), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n270), .B(KEYINPUT121), .Z(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n596), .A2(G900), .A3(G953), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT123), .B1(new_n753), .B2(new_n829), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n753), .A2(KEYINPUT123), .A3(new_n829), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n798), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n790), .A2(new_n796), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n784), .A2(new_n786), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(new_n647), .A3(new_n701), .A4(new_n741), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT124), .A4(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  INV_X1    g797(.A(new_n798), .ZN(new_n984));
  INV_X1    g798(.A(new_n977), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n975), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n790), .A2(new_n981), .A3(new_n796), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n973), .B(new_n974), .C1(new_n989), .C2(G953), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n771), .A2(new_n630), .A3(new_n681), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n500), .A3(new_n814), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT122), .Z(new_n993));
  INV_X1    g807(.A(new_n706), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n706), .B2(new_n798), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n255), .A3(new_n979), .ZN(new_n999));
  NAND3_X1  g813(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n1000), .A3(new_n972), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n990), .A2(new_n1001), .ZN(G72));
  OR2_X1    g816(.A1(new_n833), .A2(new_n841), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n685), .B(KEYINPUT63), .Z(new_n1004));
  NAND2_X1  g818(.A1(new_n412), .A2(new_n436), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT125), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n998), .A2(new_n818), .A3(new_n979), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n405), .A2(new_n411), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AND4_X1   g825(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .A4(new_n333), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n334), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1007), .B1(new_n1013), .B2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n982), .A2(new_n988), .A3(new_n818), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1011), .B(new_n333), .C1(new_n1016), .C2(new_n1004), .ZN(new_n1017));
  OAI21_X1  g831(.A(KEYINPUT126), .B1(new_n1017), .B2(new_n904), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1004), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n1010), .A3(new_n334), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1020), .A2(new_n1021), .A3(new_n943), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1006), .B(new_n1015), .C1(new_n1018), .C2(new_n1022), .ZN(G57));
endmodule


