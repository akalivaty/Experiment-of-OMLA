//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n199), .A2(new_n200), .A3(G101), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT0), .B(G128), .Z(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT70), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT70), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n207), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n201), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT78), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n194), .A2(new_n197), .A3(new_n221), .A4(new_n198), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT78), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n199), .A2(new_n223), .A3(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n203), .A3(new_n205), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n202), .A3(G143), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n204), .B(G146), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n193), .A2(G107), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n196), .A2(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n222), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n222), .A2(new_n235), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n232), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n232), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n226), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT81), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT64), .B1(new_n247), .B2(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT11), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT64), .B(new_n251), .C1(new_n247), .C2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(KEYINPUT66), .A3(new_n250), .A4(new_n252), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(G131), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT65), .B(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n249), .A2(new_n258), .A3(new_n250), .A4(new_n252), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n226), .A2(new_n241), .A3(new_n261), .A4(new_n244), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n226), .A2(new_n244), .A3(new_n241), .ZN(new_n264));
  INV_X1    g078(.A(new_n259), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n253), .B2(new_n254), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT80), .B(new_n265), .C1(new_n267), .C2(new_n256), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n257), .B2(new_n259), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n263), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n265), .B1(new_n267), .B2(new_n256), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n222), .A2(new_n235), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(new_n232), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n276), .A2(new_n230), .A3(new_n229), .A4(new_n231), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n242), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n260), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n272), .A2(new_n192), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n187), .B(new_n188), .C1(new_n273), .C2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n187), .A2(new_n188), .ZN(new_n285));
  INV_X1    g099(.A(new_n192), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n264), .B2(new_n271), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n260), .A2(KEYINPUT80), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n275), .A2(new_n269), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n275), .A2(new_n277), .A3(new_n274), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n260), .B2(new_n280), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n290), .A2(new_n245), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n263), .A2(new_n287), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n285), .B1(new_n294), .B2(G469), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT77), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT82), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT83), .Z(new_n303));
  NAND3_X1  g117(.A1(new_n296), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n232), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n203), .A2(new_n205), .B1(new_n212), .B2(new_n206), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n310));
  OAI21_X1  g124(.A(G125), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n190), .A2(G224), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n308), .B2(new_n311), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT7), .B1(new_n190), .B2(G224), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT7), .ZN(new_n317));
  AND4_X1   g131(.A1(new_n317), .A2(new_n308), .A3(new_n311), .A4(new_n312), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT69), .A2(G119), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT69), .A2(G119), .ZN(new_n321));
  OAI21_X1  g135(.A(G116), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(KEYINPUT5), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT69), .B(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G116), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(G113), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT2), .A2(G113), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(KEYINPUT2), .A2(G113), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n322), .A4(new_n324), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n334), .A3(new_n239), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT84), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n329), .A2(new_n239), .A3(new_n337), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n333), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n322), .A2(new_n324), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n201), .B1(new_n342), .B2(new_n334), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n225), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G122), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n329), .A2(new_n334), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n276), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n335), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n345), .B(KEYINPUT8), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n329), .A2(new_n239), .A3(KEYINPUT86), .A4(new_n334), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n319), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n354), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT87), .B1(new_n354), .B2(new_n188), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n339), .A2(new_n344), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n345), .B(KEYINPUT85), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n336), .A2(new_n338), .B1(new_n225), .B2(new_n343), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n359), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(new_n346), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n313), .A2(new_n314), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n306), .B1(new_n357), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n354), .A2(new_n188), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(new_n367), .A3(new_n306), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n305), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n373), .A2(KEYINPUT88), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n304), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n342), .A2(new_n334), .ZN(new_n379));
  INV_X1    g193(.A(new_n217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n216), .B1(new_n215), .B2(new_n207), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n275), .A2(new_n382), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n247), .A2(KEYINPUT67), .A3(G137), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT67), .B1(new_n247), .B2(G137), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n250), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G131), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n259), .A3(new_n232), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n379), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n379), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n388), .C1(new_n275), .C2(new_n382), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT28), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT28), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n211), .A2(new_n217), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n260), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n398), .B2(new_n388), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n396), .B(new_n388), .C1(new_n275), .C2(new_n382), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n391), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(G237), .A2(G953), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G210), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n221), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(KEYINPUT29), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n188), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n411));
  INV_X1    g225(.A(new_n210), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n257), .B2(new_n259), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n411), .B(new_n379), .C1(new_n413), .C2(new_n389), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n392), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n388), .B1(new_n275), .B2(new_n412), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n411), .B1(new_n416), .B2(new_n379), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT28), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n402), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n408), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT30), .B(new_n388), .C1(new_n275), .C2(new_n382), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n389), .B1(new_n260), .B2(new_n210), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n379), .B(new_n421), .C1(new_n422), .C2(KEYINPUT30), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n423), .A2(new_n392), .ZN(new_n424));
  INV_X1    g238(.A(new_n408), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G472), .B1(new_n410), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G472), .A2(G902), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n392), .A3(new_n408), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT31), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT31), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n423), .A2(new_n432), .A3(new_n392), .A4(new_n408), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n408), .B1(new_n418), .B2(new_n402), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT32), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT32), .B1(new_n436), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n428), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n307), .A2(G140), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT16), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G125), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(G125), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT75), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n202), .B(new_n443), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(G146), .B1(new_n453), .B2(new_n442), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n326), .A2(G128), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n227), .A2(G119), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT24), .B(G110), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(KEYINPUT23), .A3(new_n457), .ZN(new_n461));
  OR3_X1    g275(.A1(new_n326), .A2(KEYINPUT23), .A3(G128), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(G110), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n441), .A2(new_n446), .A3(G146), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G110), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n458), .A2(new_n459), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n454), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G137), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n464), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n464), .B2(new_n469), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT25), .B1(new_n476), .B2(G902), .ZN(new_n477));
  NAND2_X1  g291(.A1(G217), .A2(G902), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(G234), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT74), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n188), .C1(new_n474), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n482), .A2(G902), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n474), .B2(new_n475), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G475), .ZN(new_n490));
  INV_X1    g304(.A(new_n258), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n404), .A2(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT90), .A2(G143), .ZN(new_n493));
  OR2_X1    g307(.A1(KEYINPUT90), .A2(G143), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n493), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G214), .A3(new_n404), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n258), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT17), .B(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n503), .A2(new_n452), .A3(new_n454), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n193), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n466), .B1(new_n450), .B2(new_n202), .ZN(new_n508));
  AND4_X1   g322(.A1(KEYINPUT18), .A2(new_n500), .A3(G131), .A4(new_n501), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n500), .A2(new_n501), .B1(KEYINPUT18), .B2(G131), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n497), .A2(new_n502), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n441), .A2(new_n446), .A3(KEYINPUT19), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n450), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n513), .B(new_n454), .C1(new_n516), .C2(G146), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n507), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n490), .B(new_n188), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(KEYINPUT20), .B2(new_n519), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n507), .B1(new_n505), .B2(new_n511), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n188), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G475), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n204), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n227), .A2(G143), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G128), .B(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT91), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n534), .A3(new_n247), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT91), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT91), .B1(new_n528), .B2(new_n529), .ZN(new_n537));
  OAI21_X1  g351(.A(G134), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n323), .A2(G122), .ZN(new_n540));
  INV_X1    g354(.A(G122), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G116), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n196), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT14), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n323), .B2(G122), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n542), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(G116), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT92), .B(new_n550), .C1(new_n542), .C2(new_n546), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n539), .B(new_n544), .C1(new_n196), .C2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n543), .B(new_n196), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n533), .A2(KEYINPUT13), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(G134), .C1(KEYINPUT13), .C2(new_n528), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n535), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n297), .A2(new_n479), .A3(G953), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n557), .A3(new_n559), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(KEYINPUT93), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n553), .A2(new_n564), .A3(new_n557), .A4(new_n559), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n188), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT94), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  INV_X1    g385(.A(new_n569), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n566), .A2(new_n567), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n190), .A2(G952), .ZN(new_n577));
  NAND2_X1  g391(.A1(G234), .A2(G237), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT21), .B(G898), .Z(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(G902), .A3(G953), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n527), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n378), .A2(new_n440), .A3(new_n489), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n563), .A2(new_n586), .A3(new_n565), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n561), .A2(KEYINPUT33), .A3(new_n562), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(G478), .A3(new_n188), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n566), .A2(new_n568), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n526), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT96), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n597), .A3(new_n526), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n582), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n188), .B1(new_n434), .B2(new_n435), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(new_n436), .ZN(new_n603));
  INV_X1    g417(.A(new_n302), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n368), .B2(new_n374), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n296), .A2(new_n300), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n600), .A2(new_n489), .A3(new_n603), .A4(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  XNOR2_X1  g424(.A(new_n582), .B(KEYINPUT98), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND4_X1   g426(.A1(new_n436), .A2(new_n602), .A3(new_n489), .A4(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n553), .A2(new_n557), .A3(new_n559), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n559), .B1(new_n553), .B2(new_n557), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n614), .A2(new_n615), .A3(new_n564), .ZN(new_n616));
  INV_X1    g430(.A(new_n565), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n618), .A2(KEYINPUT94), .A3(new_n188), .A4(new_n572), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n569), .B1(new_n566), .B2(new_n567), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n574), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(new_n525), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n517), .A2(new_n511), .ZN(new_n623));
  INV_X1    g437(.A(new_n507), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n520), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n490), .A3(new_n188), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n521), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  OR3_X1    g445(.A1(new_n519), .A2(new_n630), .A3(new_n520), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n613), .A2(new_n607), .A3(new_n622), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n464), .A2(new_n469), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n486), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n485), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n378), .A2(new_n583), .A3(new_n603), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  XNOR2_X1  g459(.A(new_n579), .B(KEYINPUT100), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(G900), .B2(new_n581), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n633), .A2(new_n621), .A3(new_n525), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT101), .Z(new_n650));
  NAND3_X1  g464(.A1(new_n440), .A2(new_n607), .A3(new_n642), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n227), .ZN(G30));
  NAND3_X1  g467(.A1(new_n371), .A2(new_n367), .A3(new_n372), .ZN(new_n654));
  INV_X1    g468(.A(new_n306), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT88), .B1(new_n656), .B2(new_n373), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n376), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n302), .A3(new_n642), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n299), .B1(new_n284), .B2(new_n295), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n648), .B(KEYINPUT39), .Z(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT40), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n436), .A2(new_n437), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT32), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT32), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n424), .A2(new_n425), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n188), .B1(new_n393), .B2(new_n408), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n527), .A2(new_n576), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n660), .A2(new_n665), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  AND3_X1   g491(.A1(new_n594), .A2(new_n526), .A3(new_n648), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n440), .A2(new_n607), .A3(new_n678), .A4(new_n642), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  OAI21_X1  g494(.A(new_n188), .B1(new_n273), .B2(new_n283), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n300), .A3(new_n284), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n605), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n440), .A2(new_n684), .A3(new_n489), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n599), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT41), .B(G113), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  AOI21_X1  g502(.A(new_n488), .B1(new_n670), .B2(new_n428), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n622), .A2(new_n633), .A3(new_n612), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(KEYINPUT102), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n440), .A2(new_n684), .A3(new_n690), .A4(new_n489), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT103), .B(G116), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G18));
  NAND4_X1  g511(.A1(new_n440), .A2(new_n684), .A3(new_n583), .A4(new_n642), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND2_X1  g513(.A1(new_n656), .A2(new_n373), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n700), .A2(new_n604), .A3(new_n621), .A4(new_n526), .ZN(new_n701));
  INV_X1    g515(.A(new_n683), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n403), .A2(new_n408), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n429), .B1(new_n703), .B2(new_n434), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n602), .A2(new_n489), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n701), .A2(new_n612), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND2_X1  g521(.A1(new_n602), .A2(new_n704), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n684), .A2(new_n678), .A3(new_n642), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  XNOR2_X1  g525(.A(new_n436), .B(KEYINPUT32), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n488), .B1(new_n712), .B2(new_n428), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n657), .A2(new_n606), .A3(new_n376), .A4(new_n302), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT42), .A4(new_n678), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n440), .A3(new_n489), .A4(new_n678), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  XNOR2_X1  g536(.A(new_n649), .B(KEYINPUT101), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n714), .A3(new_n440), .A4(new_n489), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  NOR3_X1   g539(.A1(new_n657), .A2(new_n376), .A3(new_n302), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n594), .A2(new_n527), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT43), .ZN(new_n729));
  INV_X1    g543(.A(new_n603), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n642), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  OR3_X1    g546(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT106), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n732), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n294), .B(KEYINPUT45), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  INV_X1    g552(.A(new_n285), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n284), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n300), .A3(new_n663), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n735), .A2(new_n736), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n300), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n594), .A2(new_n526), .A3(new_n648), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n727), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n670), .A3(new_n428), .A4(new_n488), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  NAND2_X1  g569(.A1(new_n682), .A2(new_n284), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n728), .B1(new_n756), .B2(KEYINPUT49), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(KEYINPUT49), .ZN(new_n758));
  INV_X1    g572(.A(new_n303), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n757), .A2(new_n758), .A3(new_n488), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n674), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n300), .A3(new_n761), .A4(new_n659), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n727), .A2(new_n683), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OR4_X1    g578(.A1(new_n488), .A2(new_n764), .A3(new_n579), .A4(new_n674), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n526), .A3(new_n594), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n729), .A2(new_n646), .A3(new_n705), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n302), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n659), .A2(new_n702), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT113), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT50), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT113), .B(new_n772), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n729), .A2(new_n763), .A3(new_n646), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT114), .Z(new_n776));
  INV_X1    g590(.A(new_n642), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n776), .A2(new_n777), .A3(new_n708), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n750), .A2(new_n751), .B1(new_n300), .B2(new_n756), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n726), .A3(new_n767), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n774), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n778), .A4(new_n780), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(new_n577), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n765), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n596), .A3(new_n598), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n767), .A2(new_n684), .ZN(new_n788));
  INV_X1    g602(.A(new_n713), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n776), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT48), .Z(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n787), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n698), .B(new_n706), .C1(new_n685), .C2(new_n599), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n694), .B2(new_n691), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n621), .A2(new_n522), .A3(new_n525), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n595), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n378), .A2(new_n613), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n724), .A2(new_n584), .A3(new_n643), .A4(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n631), .A2(new_n632), .A3(new_n525), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n576), .A3(KEYINPUT107), .A4(new_n648), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT107), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n619), .B(new_n648), .C1(new_n620), .C2(new_n574), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n631), .A2(new_n632), .A3(new_n525), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n806), .A2(new_n440), .B1(new_n678), .B2(new_n709), .ZN(new_n807));
  INV_X1    g621(.A(new_n714), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n777), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n721), .A2(new_n795), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n721), .A2(KEYINPUT108), .A3(new_n795), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n679), .B(new_n710), .C1(new_n650), .C2(new_n651), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n777), .A2(new_n661), .A3(new_n648), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n605), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n777), .A2(new_n661), .A3(new_n648), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT109), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n674), .A3(new_n675), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n777), .B1(new_n670), .B2(new_n428), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n607), .C1(new_n723), .C2(new_n678), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n710), .A4(new_n822), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n815), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n829), .B1(new_n813), .B2(new_n814), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n793), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT110), .B1(new_n799), .B2(new_n809), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n721), .A2(new_n837), .A3(KEYINPUT53), .A4(new_n795), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n584), .A2(new_n643), .A3(new_n798), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n801), .A2(new_n805), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n670), .B2(new_n428), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n752), .A2(new_n708), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n642), .B(new_n714), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n839), .A2(new_n840), .A3(new_n844), .A4(new_n724), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n824), .A3(new_n828), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT111), .B1(new_n838), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n845), .A2(new_n824), .A3(new_n828), .ZN(new_n848));
  INV_X1    g662(.A(new_n794), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n695), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n716), .A2(new_n718), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT104), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n854), .B2(new_n715), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT111), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n839), .A2(new_n724), .A3(new_n844), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n832), .B1(new_n857), .B2(KEYINPUT110), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n848), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n793), .C1(new_n834), .C2(KEYINPUT53), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT112), .B1(new_n836), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n861), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n792), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n762), .B1(new_n869), .B2(new_n870), .ZN(G75));
  AOI21_X1  g685(.A(new_n188), .B1(new_n833), .B2(new_n860), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n365), .B(new_n366), .Z(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n190), .A2(G952), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G51));
  NAND2_X1  g694(.A1(new_n833), .A2(new_n860), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n861), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n739), .A2(KEYINPUT57), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n739), .A2(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n273), .B2(new_n283), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n872), .A2(G469), .A3(new_n737), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  INV_X1    g704(.A(new_n627), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n879), .ZN(G60));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT59), .Z(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n863), .A2(new_n868), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n587), .A2(new_n588), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n883), .A2(new_n587), .A3(new_n588), .A4(new_n897), .ZN(new_n903));
  INV_X1    g717(.A(new_n879), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(G63));
  XOR2_X1   g720(.A(new_n478), .B(KEYINPUT60), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n881), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n476), .B(KEYINPUT118), .Z(new_n909));
  AOI21_X1  g723(.A(new_n879), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n640), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n640), .A2(new_n911), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n881), .A2(new_n912), .A3(new_n907), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT116), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(G66));
  AOI21_X1  g731(.A(new_n190), .B1(new_n580), .B2(G224), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n795), .A2(new_n839), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n190), .ZN(new_n920));
  INV_X1    g734(.A(new_n365), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(G898), .B2(new_n190), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT119), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n920), .B(new_n923), .ZN(G69));
  AOI21_X1  g738(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT123), .Z(new_n926));
  OAI21_X1  g740(.A(new_n421), .B1(new_n422), .B2(KEYINPUT30), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n516), .ZN(new_n928));
  NAND2_X1  g742(.A1(G900), .A2(G953), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n754), .A2(new_n721), .A3(new_n724), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n816), .B(KEYINPUT120), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n745), .A2(new_n701), .A3(new_n713), .A4(new_n746), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n930), .A2(new_n747), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n928), .B(new_n929), .C1(new_n933), .C2(G953), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n689), .A2(new_n663), .A3(new_n714), .A4(new_n797), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n747), .A2(new_n754), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n931), .A2(new_n676), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n934), .B1(new_n944), .B2(new_n928), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n936), .B(new_n945), .Z(G72));
  AOI21_X1  g760(.A(new_n671), .B1(new_n833), .B2(new_n835), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n948));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n426), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT127), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n933), .B2(new_n919), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n426), .B(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n940), .A2(new_n942), .A3(new_n795), .A4(new_n839), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n951), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(KEYINPUT125), .A3(new_n951), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n671), .A3(new_n961), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n904), .A2(new_n953), .A3(new_n956), .A4(new_n962), .ZN(G57));
endmodule


