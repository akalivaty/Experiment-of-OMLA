

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(KEYINPUT29), .ZN(n671) );
  INV_X1 U549 ( .A(n977), .ZN(n708) );
  AND2_X1 U550 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U551 ( .A1(n627), .A2(n626), .ZN(n653) );
  NOR2_X1 U552 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U553 ( .A(KEYINPUT0), .B(G543), .Z(n581) );
  INV_X1 U554 ( .A(G2105), .ZN(n514) );
  OR2_X1 U555 ( .A1(n536), .A2(n581), .ZN(n532) );
  NOR2_X1 U556 ( .A1(G651), .A2(n581), .ZN(n772) );
  NOR2_X1 U557 ( .A1(G2104), .A2(n514), .ZN(n872) );
  XNOR2_X1 U558 ( .A(n643), .B(KEYINPUT15), .ZN(n988) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n769) );
  NOR2_X1 U560 ( .A1(n522), .A2(n521), .ZN(G160) );
  AND2_X1 U561 ( .A1(n514), .A2(G2104), .ZN(n867) );
  NAND2_X1 U562 ( .A1(G101), .A2(n867), .ZN(n513) );
  XOR2_X1 U563 ( .A(KEYINPUT23), .B(n513), .Z(n517) );
  NAND2_X1 U564 ( .A1(G125), .A2(n872), .ZN(n515) );
  XOR2_X1 U565 ( .A(KEYINPUT65), .B(n515), .Z(n516) );
  NAND2_X1 U566 ( .A1(n517), .A2(n516), .ZN(n522) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n518), .Z(n868) );
  NAND2_X1 U569 ( .A1(n868), .A2(G137), .ZN(n520) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U571 ( .A1(n873), .A2(G113), .ZN(n519) );
  NAND2_X1 U572 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n867), .A2(G102), .ZN(n523) );
  XNOR2_X1 U574 ( .A(n523), .B(KEYINPUT88), .ZN(n525) );
  NAND2_X1 U575 ( .A1(G138), .A2(n868), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G126), .A2(n872), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G114), .A2(n873), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U580 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U581 ( .A1(G86), .A2(n769), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G48), .A2(n772), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n535) );
  INV_X1 U584 ( .A(G651), .ZN(n536) );
  XOR2_X1 U585 ( .A(KEYINPUT66), .B(n532), .Z(n773) );
  NAND2_X1 U586 ( .A1(n773), .A2(G73), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT2), .B(n533), .Z(n534) );
  NOR2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(n536), .ZN(n538) );
  XNOR2_X1 U590 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n538), .B(n537), .ZN(n768) );
  NAND2_X1 U592 ( .A1(n768), .A2(G61), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(G305) );
  NAND2_X1 U594 ( .A1(G53), .A2(n772), .ZN(n541) );
  XOR2_X1 U595 ( .A(KEYINPUT70), .B(n541), .Z(n546) );
  NAND2_X1 U596 ( .A1(G91), .A2(n769), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G78), .A2(n773), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT69), .B(n544), .Z(n545) );
  NOR2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n768), .A2(G65), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U603 ( .A1(n769), .A2(G90), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n549), .B(KEYINPUT68), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G77), .A2(n773), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT9), .B(n552), .ZN(n556) );
  NAND2_X1 U608 ( .A1(G64), .A2(n768), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G52), .A2(n772), .ZN(n553) );
  AND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(G301) );
  INV_X1 U612 ( .A(G301), .ZN(G171) );
  XOR2_X1 U613 ( .A(KEYINPUT4), .B(KEYINPUT72), .Z(n558) );
  NAND2_X1 U614 ( .A1(G89), .A2(n769), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G76), .A2(n773), .ZN(n559) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(n559), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(KEYINPUT74), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n563), .B(n562), .ZN(n570) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(KEYINPUT76), .Z(n568) );
  NAND2_X1 U622 ( .A1(n772), .A2(G51), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT75), .B(n564), .Z(n566) );
  NAND2_X1 U624 ( .A1(n768), .A2(G63), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U626 ( .A(n568), .B(n567), .Z(n569) );
  NOR2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n571), .B(KEYINPUT77), .ZN(n572) );
  XNOR2_X1 U629 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G62), .A2(n768), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G50), .A2(n772), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U634 ( .A(KEYINPUT82), .B(n575), .ZN(n578) );
  NAND2_X1 U635 ( .A1(G75), .A2(n773), .ZN(n576) );
  XNOR2_X1 U636 ( .A(KEYINPUT83), .B(n576), .ZN(n577) );
  NOR2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n769), .A2(G88), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(G303) );
  NAND2_X1 U640 ( .A1(G49), .A2(n772), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G87), .A2(n581), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U643 ( .A1(n768), .A2(n584), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT81), .B(n585), .Z(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G288) );
  AND2_X1 U647 ( .A1(n768), .A2(G60), .ZN(n591) );
  NAND2_X1 U648 ( .A1(G85), .A2(n769), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G47), .A2(n772), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U651 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G72), .A2(n773), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n627) );
  NOR2_X1 U655 ( .A1(G1384), .A2(G164), .ZN(n594) );
  XNOR2_X1 U656 ( .A(n594), .B(KEYINPUT64), .ZN(n625) );
  NOR2_X1 U657 ( .A1(n627), .A2(n625), .ZN(n739) );
  NAND2_X1 U658 ( .A1(G104), .A2(n867), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G140), .A2(n868), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U661 ( .A(KEYINPUT34), .B(n597), .ZN(n602) );
  NAND2_X1 U662 ( .A1(G128), .A2(n872), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G116), .A2(n873), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U665 ( .A(KEYINPUT35), .B(n600), .Z(n601) );
  NOR2_X1 U666 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U667 ( .A(KEYINPUT36), .B(n603), .ZN(n883) );
  XOR2_X1 U668 ( .A(G2067), .B(KEYINPUT37), .Z(n604) );
  XNOR2_X1 U669 ( .A(KEYINPUT89), .B(n604), .ZN(n737) );
  NOR2_X1 U670 ( .A1(n883), .A2(n737), .ZN(n949) );
  NAND2_X1 U671 ( .A1(n739), .A2(n949), .ZN(n735) );
  NAND2_X1 U672 ( .A1(G119), .A2(n872), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G107), .A2(n873), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n868), .A2(G131), .ZN(n607) );
  XOR2_X1 U676 ( .A(KEYINPUT90), .B(n607), .Z(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n867), .A2(G95), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n862) );
  NAND2_X1 U680 ( .A1(G1991), .A2(n862), .ZN(n621) );
  NAND2_X1 U681 ( .A1(G105), .A2(n867), .ZN(n612) );
  XOR2_X1 U682 ( .A(KEYINPUT38), .B(n612), .Z(n617) );
  NAND2_X1 U683 ( .A1(G129), .A2(n872), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G117), .A2(n873), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT91), .B(n615), .Z(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n868), .A2(G141), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n858) );
  NAND2_X1 U690 ( .A1(G1996), .A2(n858), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT92), .B(n622), .Z(n953) );
  XNOR2_X1 U693 ( .A(KEYINPUT93), .B(n739), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n953), .A2(n623), .ZN(n731) );
  INV_X1 U695 ( .A(n731), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n735), .A2(n624), .ZN(n726) );
  INV_X1 U697 ( .A(n625), .ZN(n626) );
  INV_X1 U698 ( .A(n653), .ZN(n694) );
  NAND2_X1 U699 ( .A1(G8), .A2(n694), .ZN(n719) );
  NOR2_X1 U700 ( .A1(G1981), .A2(G305), .ZN(n628) );
  XOR2_X1 U701 ( .A(n628), .B(KEYINPUT24), .Z(n629) );
  NOR2_X1 U702 ( .A1(n719), .A2(n629), .ZN(n724) );
  NOR2_X1 U703 ( .A1(G2084), .A2(n694), .ZN(n678) );
  NAND2_X1 U704 ( .A1(G8), .A2(n678), .ZN(n692) );
  NOR2_X1 U705 ( .A1(G1966), .A2(n719), .ZN(n690) );
  INV_X1 U706 ( .A(G299), .ZN(n985) );
  NAND2_X1 U707 ( .A1(n653), .A2(G2072), .ZN(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT27), .B(n630), .Z(n632) );
  NAND2_X1 U709 ( .A1(n694), .A2(G1956), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT95), .ZN(n635) );
  OR2_X1 U712 ( .A1(n985), .A2(n635), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n634), .B(KEYINPUT28), .ZN(n670) );
  NAND2_X1 U714 ( .A1(n985), .A2(n635), .ZN(n668) );
  NAND2_X1 U715 ( .A1(G54), .A2(n772), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G66), .A2(n768), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G92), .A2(n769), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n773), .A2(G79), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT71), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G56), .A2(n768), .ZN(n644) );
  XOR2_X1 U724 ( .A(KEYINPUT14), .B(n644), .Z(n650) );
  NAND2_X1 U725 ( .A1(n769), .A2(G81), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT12), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G68), .A2(n773), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U729 ( .A(KEYINPUT13), .B(n648), .Z(n649) );
  NOR2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n772), .A2(G43), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n971) );
  AND2_X1 U733 ( .A1(n653), .A2(G1996), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n694), .A2(G1341), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U738 ( .A1(n971), .A2(n658), .ZN(n659) );
  OR2_X1 U739 ( .A1(n988), .A2(n659), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n988), .A2(n659), .ZN(n664) );
  AND2_X1 U741 ( .A1(n653), .A2(G2067), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n660), .B(KEYINPUT97), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n694), .A2(G1348), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n672), .B(n671), .ZN(n677) );
  INV_X1 U750 ( .A(G1961), .ZN(n989) );
  NAND2_X1 U751 ( .A1(n694), .A2(n989), .ZN(n674) );
  XNOR2_X1 U752 ( .A(G2078), .B(KEYINPUT25), .ZN(n899) );
  NAND2_X1 U753 ( .A1(n653), .A2(n899), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n682) );
  AND2_X1 U755 ( .A1(n682), .A2(G171), .ZN(n675) );
  XOR2_X1 U756 ( .A(KEYINPUT94), .B(n675), .Z(n676) );
  NAND2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n690), .A2(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G8), .A2(n679), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT30), .B(n680), .ZN(n681) );
  NOR2_X1 U761 ( .A1(G168), .A2(n681), .ZN(n684) );
  NOR2_X1 U762 ( .A1(G171), .A2(n682), .ZN(n683) );
  NOR2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U764 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n685) );
  XNOR2_X1 U765 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n693) );
  XNOR2_X1 U767 ( .A(KEYINPUT99), .B(n693), .ZN(n689) );
  NOR2_X1 U768 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n692), .A2(n691), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n693), .A2(G286), .ZN(n699) );
  NOR2_X1 U771 ( .A1(G1971), .A2(n719), .ZN(n696) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n694), .ZN(n695) );
  NOR2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U774 ( .A1(n697), .A2(G303), .ZN(n698) );
  NAND2_X1 U775 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U776 ( .A1(n700), .A2(G8), .ZN(n701) );
  XNOR2_X1 U777 ( .A(n701), .B(KEYINPUT32), .ZN(n702) );
  NAND2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n718) );
  NOR2_X1 U779 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NOR2_X1 U780 ( .A1(G1971), .A2(G303), .ZN(n704) );
  NOR2_X1 U781 ( .A1(n972), .A2(n704), .ZN(n705) );
  XNOR2_X1 U782 ( .A(KEYINPUT100), .B(n705), .ZN(n706) );
  NAND2_X1 U783 ( .A1(n718), .A2(n706), .ZN(n710) );
  NAND2_X1 U784 ( .A1(G288), .A2(G1976), .ZN(n707) );
  XOR2_X1 U785 ( .A(KEYINPUT101), .B(n707), .Z(n977) );
  NOR2_X1 U786 ( .A1(n719), .A2(n708), .ZN(n709) );
  NOR2_X1 U787 ( .A1(KEYINPUT33), .A2(n711), .ZN(n714) );
  NAND2_X1 U788 ( .A1(n972), .A2(KEYINPUT33), .ZN(n712) );
  NOR2_X1 U789 ( .A1(n712), .A2(n719), .ZN(n713) );
  NOR2_X1 U790 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U791 ( .A(G1981), .B(G305), .Z(n981) );
  NAND2_X1 U792 ( .A1(n715), .A2(n981), .ZN(n722) );
  NOR2_X1 U793 ( .A1(G2090), .A2(G303), .ZN(n716) );
  NAND2_X1 U794 ( .A1(G8), .A2(n716), .ZN(n717) );
  NAND2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U798 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U799 ( .A(G1986), .B(G290), .ZN(n976) );
  NAND2_X1 U800 ( .A1(n976), .A2(n739), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n742) );
  NOR2_X1 U802 ( .A1(G1991), .A2(n862), .ZN(n948) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n729) );
  NOR2_X1 U804 ( .A1(n948), .A2(n729), .ZN(n730) );
  NOR2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n858), .ZN(n962) );
  NOR2_X1 U807 ( .A1(n732), .A2(n962), .ZN(n733) );
  XNOR2_X1 U808 ( .A(n733), .B(KEYINPUT39), .ZN(n734) );
  XNOR2_X1 U809 ( .A(n734), .B(KEYINPUT102), .ZN(n736) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U811 ( .A1(n883), .A2(n737), .ZN(n954) );
  NAND2_X1 U812 ( .A1(n738), .A2(n954), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U816 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U817 ( .A(G57), .ZN(G237) );
  INV_X1 U818 ( .A(G132), .ZN(G219) );
  INV_X1 U819 ( .A(G82), .ZN(G220) );
  NAND2_X1 U820 ( .A1(G7), .A2(G661), .ZN(n744) );
  XNOR2_X1 U821 ( .A(n744), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U822 ( .A(G223), .ZN(n816) );
  NAND2_X1 U823 ( .A1(n816), .A2(G567), .ZN(n745) );
  XOR2_X1 U824 ( .A(KEYINPUT11), .B(n745), .Z(G234) );
  INV_X1 U825 ( .A(G860), .ZN(n750) );
  OR2_X1 U826 ( .A1(n971), .A2(n750), .ZN(G153) );
  NAND2_X1 U827 ( .A1(G868), .A2(G301), .ZN(n747) );
  OR2_X1 U828 ( .A1(n988), .A2(G868), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n747), .A2(n746), .ZN(G284) );
  INV_X1 U830 ( .A(G868), .ZN(n789) );
  NOR2_X1 U831 ( .A1(G286), .A2(n789), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G868), .A2(G299), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n749), .A2(n748), .ZN(G297) );
  NAND2_X1 U834 ( .A1(n750), .A2(G559), .ZN(n751) );
  NAND2_X1 U835 ( .A1(n751), .A2(n988), .ZN(n752) );
  XNOR2_X1 U836 ( .A(n752), .B(KEYINPUT78), .ZN(n753) );
  XNOR2_X1 U837 ( .A(KEYINPUT16), .B(n753), .ZN(G148) );
  NOR2_X1 U838 ( .A1(G868), .A2(n971), .ZN(n756) );
  NAND2_X1 U839 ( .A1(n988), .A2(G868), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G559), .A2(n754), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n756), .A2(n755), .ZN(G282) );
  XOR2_X1 U842 ( .A(G2100), .B(KEYINPUT80), .Z(n766) );
  NAND2_X1 U843 ( .A1(G99), .A2(n867), .ZN(n758) );
  NAND2_X1 U844 ( .A1(G111), .A2(n873), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT79), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G135), .A2(n868), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n872), .A2(G123), .ZN(n762) );
  XOR2_X1 U850 ( .A(KEYINPUT18), .B(n762), .Z(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n947) );
  XNOR2_X1 U852 ( .A(G2096), .B(n947), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(G156) );
  NAND2_X1 U854 ( .A1(n988), .A2(G559), .ZN(n786) );
  XNOR2_X1 U855 ( .A(n971), .B(n786), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n767), .A2(G860), .ZN(n778) );
  NAND2_X1 U857 ( .A1(G67), .A2(n768), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G93), .A2(n769), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n777) );
  NAND2_X1 U860 ( .A1(n772), .A2(G55), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G80), .A2(n773), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n788) );
  XOR2_X1 U864 ( .A(n778), .B(n788), .Z(G145) );
  INV_X1 U865 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U866 ( .A(KEYINPUT19), .B(G305), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(G288), .ZN(n780) );
  XOR2_X1 U868 ( .A(n780), .B(n788), .Z(n782) );
  XNOR2_X1 U869 ( .A(G290), .B(G166), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U871 ( .A(n783), .B(G299), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(n971), .ZN(n886) );
  XOR2_X1 U873 ( .A(n886), .B(KEYINPUT84), .Z(n785) );
  XNOR2_X1 U874 ( .A(n786), .B(n785), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n787), .A2(G868), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(G295) );
  NAND2_X1 U878 ( .A1(G2084), .A2(G2078), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT20), .B(n792), .Z(n793) );
  NAND2_X1 U880 ( .A1(G2090), .A2(n793), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n794) );
  XNOR2_X1 U882 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G2072), .A2(n796), .ZN(G158) );
  XNOR2_X1 U884 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U885 ( .A1(G220), .A2(G219), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT22), .B(n797), .Z(n798) );
  NOR2_X1 U887 ( .A1(G218), .A2(n798), .ZN(n799) );
  XNOR2_X1 U888 ( .A(KEYINPUT86), .B(n799), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n800), .A2(G96), .ZN(n820) );
  NAND2_X1 U890 ( .A1(n820), .A2(G2106), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G69), .A2(G120), .ZN(n801) );
  NOR2_X1 U892 ( .A1(G237), .A2(n801), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G108), .A2(n802), .ZN(n821) );
  NAND2_X1 U894 ( .A1(n821), .A2(G567), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n822) );
  NAND2_X1 U896 ( .A1(G661), .A2(G483), .ZN(n805) );
  XOR2_X1 U897 ( .A(KEYINPUT87), .B(n805), .Z(n806) );
  NOR2_X1 U898 ( .A1(n822), .A2(n806), .ZN(n819) );
  NAND2_X1 U899 ( .A1(n819), .A2(G36), .ZN(G176) );
  XNOR2_X1 U900 ( .A(G1341), .B(G2454), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(G2430), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(G1348), .ZN(n814) );
  XOR2_X1 U903 ( .A(G2443), .B(G2427), .Z(n810) );
  XNOR2_X1 U904 ( .A(G2438), .B(G2446), .ZN(n809) );
  XNOR2_X1 U905 ( .A(n810), .B(n809), .ZN(n812) );
  XOR2_X1 U906 ( .A(G2451), .B(G2435), .Z(n811) );
  XNOR2_X1 U907 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(G14), .ZN(n891) );
  XNOR2_X1 U910 ( .A(KEYINPUT103), .B(n891), .ZN(G401) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U913 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  INV_X1 U922 ( .A(n822), .ZN(G319) );
  XNOR2_X1 U923 ( .A(G1981), .B(KEYINPUT41), .ZN(n832) );
  XOR2_X1 U924 ( .A(G1976), .B(G1971), .Z(n824) );
  XNOR2_X1 U925 ( .A(G1986), .B(G1956), .ZN(n823) );
  XNOR2_X1 U926 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U927 ( .A(G1961), .B(G1966), .Z(n826) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1991), .ZN(n825) );
  XNOR2_X1 U929 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U930 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U931 ( .A(KEYINPUT106), .B(G2474), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(G229) );
  XOR2_X1 U934 ( .A(KEYINPUT104), .B(G2678), .Z(n834) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n833) );
  XNOR2_X1 U936 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(G2090), .Z(n836) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U940 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2100), .B(G2096), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U943 ( .A(G2084), .B(G2078), .Z(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(G227) );
  NAND2_X1 U945 ( .A1(G124), .A2(n872), .ZN(n843) );
  XOR2_X1 U946 ( .A(KEYINPUT44), .B(n843), .Z(n844) );
  XNOR2_X1 U947 ( .A(n844), .B(KEYINPUT107), .ZN(n846) );
  NAND2_X1 U948 ( .A1(G100), .A2(n867), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G112), .A2(n873), .ZN(n848) );
  NAND2_X1 U951 ( .A1(G136), .A2(n868), .ZN(n847) );
  NAND2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U953 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U954 ( .A1(G130), .A2(n872), .ZN(n852) );
  NAND2_X1 U955 ( .A1(G118), .A2(n873), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G106), .A2(n867), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G142), .A2(n868), .ZN(n853) );
  NAND2_X1 U959 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U960 ( .A(n855), .B(KEYINPUT45), .Z(n856) );
  NOR2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n947), .B(n860), .ZN(n882) );
  XOR2_X1 U964 ( .A(KEYINPUT108), .B(KEYINPUT110), .Z(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(n863), .B(KEYINPUT48), .Z(n865) );
  XNOR2_X1 U967 ( .A(G164), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(n866), .B(G162), .Z(n880) );
  NAND2_X1 U970 ( .A1(G103), .A2(n867), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G139), .A2(n868), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT109), .B(n871), .Z(n878) );
  NAND2_X1 U974 ( .A1(G127), .A2(n872), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G115), .A2(n873), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n957) );
  XNOR2_X1 U979 ( .A(G160), .B(n957), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U983 ( .A1(G37), .A2(n885), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n988), .B(G286), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(G301), .B(n888), .Z(n889) );
  NOR2_X1 U987 ( .A1(G37), .A2(n889), .ZN(n890) );
  XOR2_X1 U988 ( .A(KEYINPUT111), .B(n890), .Z(G397) );
  NAND2_X1 U989 ( .A1(G319), .A2(n891), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G229), .A2(G227), .ZN(n892) );
  XNOR2_X1 U991 ( .A(KEYINPUT49), .B(n892), .ZN(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G395), .A2(G397), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(G225) );
  INV_X1 U995 ( .A(G225), .ZN(G308) );
  INV_X1 U996 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U997 ( .A(KEYINPUT115), .B(G1996), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n897), .B(G32), .ZN(n907) );
  XOR2_X1 U999 ( .A(G2072), .B(G33), .Z(n898) );
  NAND2_X1 U1000 ( .A1(n898), .A2(G28), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(G27), .B(n899), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G26), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(G1991), .B(G25), .ZN(n900) );
  NOR2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  NOR2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(KEYINPUT53), .B(n908), .ZN(n912) );
  XOR2_X1 U1009 ( .A(G34), .B(KEYINPUT116), .Z(n910) );
  XNOR2_X1 U1010 ( .A(G2084), .B(KEYINPUT54), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT114), .B(G2090), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(G35), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1016 ( .A(KEYINPUT117), .B(n916), .Z(n917) );
  NOR2_X1 U1017 ( .A1(G29), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(KEYINPUT55), .B(n918), .ZN(n1005) );
  XOR2_X1 U1019 ( .A(G16), .B(KEYINPUT122), .Z(n944) );
  XOR2_X1 U1020 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n919) );
  XNOR2_X1 U1021 ( .A(KEYINPUT61), .B(n919), .ZN(n942) );
  XNOR2_X1 U1022 ( .A(G1348), .B(KEYINPUT59), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(n920), .B(G4), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1956), .B(G20), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(G1981), .B(G6), .ZN(n921) );
  NOR2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1028 ( .A(KEYINPUT123), .B(G1341), .Z(n925) );
  XNOR2_X1 U1029 ( .A(G19), .B(n925), .ZN(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(KEYINPUT60), .B(n928), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G1966), .B(KEYINPUT124), .ZN(n929) );
  XNOR2_X1 U1033 ( .A(n929), .B(G21), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n931) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n930) );
  NOR2_X1 U1036 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n932) );
  NAND2_X1 U1038 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1040 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(G5), .B(G1961), .ZN(n939) );
  NOR2_X1 U1043 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1044 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n945), .ZN(n1003) );
  XOR2_X1 U1047 ( .A(G2084), .B(G160), .Z(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(KEYINPUT112), .B(n952), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n968) );
  XOR2_X1 U1054 ( .A(G2072), .B(n957), .Z(n959) );
  XOR2_X1 U1055 ( .A(G164), .B(G2078), .Z(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1057 ( .A(KEYINPUT50), .B(n960), .Z(n966) );
  XOR2_X1 U1058 ( .A(G2090), .B(G162), .Z(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1060 ( .A(KEYINPUT51), .B(n963), .Z(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT113), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT52), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(G29), .ZN(n1001) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XOR2_X1 U1067 ( .A(n971), .B(G1341), .Z(n974) );
  XNOR2_X1 U1068 ( .A(n972), .B(KEYINPUT121), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT118), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n982), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n997) );
  XNOR2_X1 U1077 ( .A(G166), .B(G1971), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n985), .B(G1956), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G1348), .B(n988), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G171), .B(KEYINPUT119), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n990), .B(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT120), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(n1006), .B(KEYINPUT127), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(KEYINPUT62), .B(n1007), .ZN(G311) );
  INV_X1 U1093 ( .A(G311), .ZN(G150) );
endmodule

