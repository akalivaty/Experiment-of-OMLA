//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT86), .Z(new_n205));
  XOR2_X1   g004(.A(KEYINPUT87), .B(G22gat), .Z(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n211), .C1(new_n212), .C2(KEYINPUT2), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n208), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G211gat), .B(G218gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT72), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(G197gat), .ZN(new_n226));
  INV_X1    g025(.A(G204gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n224), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n222), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n221), .A3(new_n234), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n231), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n207), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n207), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n213), .A2(new_n221), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n228), .A2(new_n229), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n241), .A2(new_n225), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n224), .B(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT29), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n206), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n246), .A3(new_n206), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n205), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n204), .ZN(new_n251));
  INV_X1    g050(.A(G22gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n238), .B2(new_n246), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT73), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n258), .A2(G169gat), .A3(G176gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT23), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n267), .A2(new_n268), .A3(new_n271), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n260), .B1(KEYINPUT23), .B2(new_n262), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n279), .A2(new_n277), .A3(new_n259), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n271), .A2(new_n265), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n273), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT67), .B1(new_n289), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n273), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT26), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n262), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n297), .B(new_n269), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(new_n272), .B2(KEYINPUT27), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n288), .A3(G183gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n283), .A2(KEYINPUT27), .A3(new_n284), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n278), .A2(new_n287), .B1(new_n294), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n257), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n278), .A2(new_n287), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n288), .A2(G183gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT67), .ZN(new_n317));
  AOI21_X1  g116(.A(G190gat), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n308), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g119(.A(new_n311), .B(new_n257), .C1(new_n312), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n317), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n322), .B2(new_n273), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n261), .A2(new_n298), .A3(new_n262), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n297), .A2(new_n269), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n327), .A2(new_n282), .A3(new_n288), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n260), .A2(KEYINPUT23), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n258), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI211_X1 g130(.A(KEYINPUT25), .B(new_n330), .C1(new_n331), .C2(new_n260), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n285), .B2(new_n281), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT25), .B1(new_n264), .B2(new_n275), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n323), .A2(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n257), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT74), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n310), .B1(new_n321), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n243), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n329), .B1(KEYINPUT28), .B2(new_n293), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n276), .A2(new_n277), .B1(new_n280), .B2(new_n286), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n310), .A2(new_n340), .A3(new_n231), .A4(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n312), .B2(new_n320), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n231), .B(new_n343), .C1(new_n345), .C2(new_n336), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND4_X1  g149(.A1(new_n339), .A2(new_n344), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n347), .A2(new_n344), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n339), .A4(new_n350), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n344), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n311), .B1(new_n309), .B2(new_n257), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n335), .A2(KEYINPUT74), .A3(new_n336), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n231), .B1(new_n362), .B2(new_n310), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n339), .A2(KEYINPUT76), .A3(new_n344), .A4(new_n347), .ZN(new_n365));
  INV_X1    g164(.A(new_n350), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n359), .A2(new_n363), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n350), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n371), .B(KEYINPUT80), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT68), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(G120gat), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT69), .B1(new_n378), .B2(G113gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n376), .A3(G120gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n379), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(G127gat), .A2(G134gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(G127gat), .A2(G134gat), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT1), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n378), .A2(G113gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n376), .A2(G120gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n383), .A2(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n222), .A2(new_n374), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n383), .A2(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n391), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT4), .B1(new_n397), .B2(new_n240), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n222), .A2(new_n399), .A3(new_n392), .A4(new_n374), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n392), .A2(KEYINPUT78), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n236), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n373), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n404), .A3(new_n240), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n222), .A2(new_n392), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n373), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT39), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(KEYINPUT88), .A3(KEYINPUT39), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT39), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n407), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT40), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n398), .A2(new_n393), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n406), .A3(new_n373), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n410), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n372), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n428), .A2(new_n406), .A3(new_n434), .A4(new_n373), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n401), .A2(new_n431), .A3(new_n373), .A4(new_n406), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT89), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n421), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(KEYINPUT89), .A3(new_n437), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n425), .A2(new_n427), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n255), .B1(new_n370), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n364), .A2(KEYINPUT37), .A3(new_n365), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n366), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n446), .A2(KEYINPUT91), .B1(new_n368), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n450), .A3(new_n366), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n439), .B1(new_n436), .B2(new_n437), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n439), .A3(new_n437), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n455), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n352), .A2(new_n355), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n310), .A2(new_n343), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n243), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n338), .A2(new_n231), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT38), .B(new_n350), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n368), .A2(new_n448), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n443), .B1(new_n452), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n309), .A2(new_n397), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  INV_X1    g272(.A(G233gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n335), .A2(new_n392), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G15gat), .B(G43gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n477), .B(KEYINPUT32), .C1(new_n479), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n476), .ZN(new_n489));
  INV_X1    g288(.A(new_n475), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI211_X1 g290(.A(KEYINPUT34), .B(new_n475), .C1(new_n472), .C2(new_n476), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n484), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT36), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n497), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(KEYINPUT36), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n494), .A2(KEYINPUT71), .A3(new_n497), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n357), .A2(new_n367), .A3(new_n369), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n458), .A2(new_n509), .A3(new_n455), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n454), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n456), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n513), .A3(KEYINPUT85), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n453), .B1(new_n459), .B2(KEYINPUT84), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n456), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n517), .B2(new_n370), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n506), .B1(new_n519), .B2(new_n255), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n496), .A2(new_n498), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n255), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n524));
  INV_X1    g323(.A(new_n249), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n247), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n526), .A2(new_n205), .B1(new_n253), .B2(new_n251), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n501), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n528), .A2(new_n461), .A3(KEYINPUT35), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n507), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n471), .A2(new_n520), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(G1gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT96), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT96), .A3(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(KEYINPUT96), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n533), .A2(new_n535), .A3(new_n540), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT93), .B(G29gat), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT14), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT14), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT92), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n544), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n550), .B1(G36gat), .B2(new_n543), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(KEYINPUT95), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n556), .B2(new_n557), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(KEYINPUT95), .A3(new_n557), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n542), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT13), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n559), .B(KEYINPUT17), .C1(new_n562), .C2(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n542), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n539), .A3(new_n541), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n577), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n578), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G197gat), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT11), .B(G169gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT12), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n573), .A2(new_n581), .A3(new_n588), .A4(new_n582), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n531), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT97), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n595), .B(new_n596), .C1(new_n600), .C2(KEYINPUT9), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT97), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n539), .A2(new_n541), .B1(new_n607), .B2(KEYINPUT21), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT99), .ZN(new_n615));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  XNOR2_X1  g423(.A(G99gat), .B(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  AOI22_X1  g427(.A1(KEYINPUT8), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n624), .B2(new_n629), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n575), .B(new_n576), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n568), .A2(new_n633), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G190gat), .B(G218gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n637), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT100), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n629), .ZN(new_n646));
  INV_X1    g445(.A(new_n625), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n599), .A2(new_n602), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n604), .B1(new_n605), .B2(KEYINPUT97), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT101), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n603), .B(new_n606), .C1(new_n630), .C2(new_n631), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n655), .A3(new_n653), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n633), .A2(new_n657), .A3(new_n607), .A4(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n655), .ZN(new_n662));
  INV_X1    g461(.A(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n664), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n622), .A2(new_n645), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n594), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n517), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g478(.A(new_n536), .B1(new_n677), .B2(new_n370), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n676), .A2(new_n507), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT42), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n676), .B2(new_n505), .ZN(new_n685));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n501), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n676), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n527), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n622), .A2(new_n645), .A3(new_n672), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n594), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n693), .A2(new_n513), .A3(new_n543), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT45), .Z(new_n695));
  XOR2_X1   g494(.A(new_n672), .B(KEYINPUT102), .Z(new_n696));
  NOR3_X1   g495(.A1(new_n622), .A2(new_n593), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n531), .B2(new_n645), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n524), .A2(new_n530), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n519), .A2(new_n255), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n471), .A3(new_n505), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n645), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n698), .B1(new_n700), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n517), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n543), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n709), .B2(new_n517), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n695), .B1(new_n712), .B2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n693), .A2(G36gat), .A3(new_n507), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n709), .A2(new_n370), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n546), .ZN(G1329gat));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n709), .A2(new_n506), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n693), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n721), .A3(new_n501), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n720), .B2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI221_X1 g526(.A(new_n724), .B1(new_n719), .B2(KEYINPUT47), .C1(new_n720), .C2(new_n721), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n255), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G50gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n527), .A2(G50gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n693), .B2(KEYINPUT106), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT48), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n730), .A2(G50gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n736), .A2(new_n738), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n735), .A2(new_n739), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g542(.A(new_n622), .ZN(new_n744));
  INV_X1    g543(.A(new_n696), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n744), .A2(new_n745), .A3(new_n592), .A4(new_n705), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n704), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n517), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g549(.A(new_n747), .B(KEYINPUT108), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n507), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n751), .B2(new_n505), .ZN(new_n757));
  INV_X1    g556(.A(G71gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n758), .A3(new_n501), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g560(.A1(new_n751), .A2(new_n527), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT109), .B(G78gat), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n370), .A2(new_n442), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n527), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n451), .A3(new_n468), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT38), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n461), .A2(new_n462), .A3(new_n469), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n527), .B1(new_n514), .B2(new_n518), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(new_n773), .A3(new_n506), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n523), .A2(KEYINPUT35), .B1(new_n529), .B2(new_n507), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT110), .B(new_n705), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n622), .A2(new_n592), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT110), .B1(new_n704), .B2(new_n705), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n765), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n777), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n645), .B1(new_n701), .B2(new_n703), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(KEYINPUT110), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n531), .B2(new_n645), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(new_n627), .A3(new_n517), .A4(new_n672), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n777), .A2(new_n672), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n700), .B2(new_n708), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n513), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1336gat));
  NAND4_X1  g592(.A1(new_n787), .A2(new_n628), .A3(new_n370), .A4(new_n696), .ZN(new_n794));
  OAI21_X1  g593(.A(G92gat), .B1(new_n791), .B2(new_n507), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1337gat));
  NOR2_X1   g599(.A1(new_n673), .A2(G99gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n787), .A2(new_n501), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G99gat), .B1(new_n791), .B2(new_n505), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1338gat));
  NOR3_X1   g603(.A1(new_n745), .A2(new_n527), .A3(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n780), .B2(new_n786), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT53), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n778), .A2(new_n779), .A3(new_n765), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n783), .B2(new_n785), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n790), .B2(new_n255), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n810), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n807), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(new_n816), .A3(new_n810), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT112), .B1(new_n807), .B2(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1339gat));
  NAND4_X1  g623(.A1(new_n654), .A2(new_n656), .A3(new_n663), .A4(new_n658), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n659), .A2(new_n827), .A3(new_n660), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n669), .A4(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n669), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n592), .A2(new_n671), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n569), .A2(new_n572), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(KEYINPUT113), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n838), .B(new_n570), .C1(new_n577), .C2(new_n578), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n587), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n591), .A3(new_n672), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n705), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n671), .A3(new_n829), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n591), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n645), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n744), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n622), .A2(new_n593), .A3(new_n645), .A4(new_n673), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n513), .A2(new_n370), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n527), .A3(new_n501), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n593), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n522), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n592), .A2(new_n376), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT114), .Z(G1340gat));
  NOR3_X1   g655(.A1(new_n851), .A2(new_n378), .A3(new_n745), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n522), .A3(new_n672), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n378), .B2(new_n858), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n853), .A2(new_n744), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n622), .A2(G127gat), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n860), .A2(G127gat), .B1(new_n851), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT115), .ZN(G1342gat));
  NOR3_X1   g662(.A1(new_n853), .A2(G134gat), .A3(new_n645), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n705), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n866), .B2(new_n528), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n505), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT116), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n527), .B1(new_n846), .B2(new_n847), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n847), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n841), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n833), .A2(new_n878), .A3(new_n671), .A4(new_n829), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n592), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n705), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n744), .B1(new_n881), .B2(new_n845), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n744), .C1(new_n881), .C2(new_n845), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n527), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n873), .B1(new_n886), .B2(new_n871), .ZN(new_n887));
  OAI21_X1  g686(.A(G141gat), .B1(new_n887), .B2(new_n593), .ZN(new_n888));
  INV_X1    g687(.A(new_n869), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(G141gat), .A3(new_n593), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT58), .B1(new_n892), .B2(KEYINPUT122), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n888), .B(new_n893), .C1(KEYINPUT122), .C2(new_n892), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n845), .B1(new_n898), .B2(new_n645), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n883), .B1(new_n899), .B2(new_n622), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n847), .A3(new_n885), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n871), .B1(new_n901), .B2(new_n255), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n872), .A2(new_n871), .ZN(new_n903));
  INV_X1    g702(.A(new_n870), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT120), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n873), .C1(new_n886), .C2(new_n871), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n908), .A3(new_n592), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n892), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n895), .B1(new_n911), .B2(KEYINPUT58), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n891), .B1(new_n909), .B2(G141gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(KEYINPUT121), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n894), .B1(new_n912), .B2(new_n915), .ZN(G1344gat));
  NOR2_X1   g715(.A1(new_n216), .A2(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n906), .A2(new_n908), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n673), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT57), .B(new_n527), .C1(new_n882), .C2(new_n847), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n872), .A2(new_n871), .ZN(new_n921));
  NOR4_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n673), .A4(new_n870), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT59), .B1(new_n922), .B2(new_n216), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n890), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n216), .A3(new_n672), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n918), .B2(new_n744), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n209), .A3(new_n622), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(KEYINPUT123), .B1(new_n918), .B2(new_n645), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G162gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n645), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n505), .A2(new_n210), .A3(new_n255), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n866), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n507), .A2(new_n517), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n848), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n255), .A3(new_n521), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n592), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n528), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n593), .A2(new_n295), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n938), .B2(new_n672), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT124), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n745), .A2(new_n296), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n940), .B2(new_n945), .ZN(G1349gat));
  AOI22_X1  g745(.A1(new_n940), .A2(new_n622), .B1(new_n283), .B2(new_n284), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n622), .A2(new_n322), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g749(.A(new_n273), .B1(new_n940), .B2(new_n705), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT61), .Z(new_n952));
  NAND3_X1  g751(.A1(new_n938), .A2(new_n273), .A3(new_n705), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1351gat));
  AND2_X1   g753(.A1(new_n936), .A2(new_n505), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n872), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(new_n226), .A3(new_n592), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n955), .B(KEYINPUT126), .ZN(new_n959));
  OR3_X1    g758(.A1(new_n920), .A2(new_n921), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n593), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n227), .A3(new_n672), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n960), .B2(new_n745), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n956), .A2(new_n967), .A3(new_n622), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n960), .B2(new_n744), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AND2_X1   g772(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n705), .B1(new_n960), .B2(KEYINPUT127), .ZN(new_n975));
  OAI21_X1  g774(.A(G218gat), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(G218gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n956), .A2(new_n977), .A3(new_n705), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1355gat));
endmodule


