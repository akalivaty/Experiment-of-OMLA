//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1240,
    new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G221), .A2(G218), .A3(G219), .A4(G220), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n451), .B2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n465), .B(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n463), .A2(KEYINPUT72), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n482), .A3(new_n462), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n474), .B1(new_n483), .B2(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT4), .A4(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n476), .A2(new_n478), .A3(G138), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n462), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n476), .A2(new_n478), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n491), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n502), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n501), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT73), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(G543), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT74), .B1(new_n510), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(new_n515), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n518), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n505), .A2(new_n506), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n512), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  INV_X1    g110(.A(G77), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(new_n501), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n539), .B1(new_n536), .B2(new_n501), .C1(new_n534), .C2(new_n535), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(G651), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n518), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n525), .A2(G90), .B1(G52), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n500), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(G43), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n525), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND3_X1  g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n511), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n500), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n515), .A2(KEYINPUT78), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n507), .A2(new_n569), .A3(new_n511), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT79), .B1(new_n571), .B2(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n573), .B(new_n574), .C1(new_n568), .C2(new_n570), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n567), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  AND4_X1   g152(.A1(new_n569), .A2(new_n533), .A3(new_n512), .A4(new_n511), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n569), .B1(new_n507), .B2(new_n511), .ZN(new_n579));
  OAI21_X1  g154(.A(G91), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(new_n573), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n571), .A2(KEYINPUT79), .A3(G91), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(new_n584), .A3(new_n567), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(new_n585), .ZN(G299));
  OR2_X1    g161(.A1(new_n526), .A2(new_n531), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  OAI21_X1  g163(.A(G87), .B1(new_n578), .B2(new_n579), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n507), .A2(G74), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G49), .B2(new_n542), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n593), .B(G87), .C1(new_n578), .C2(new_n579), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n534), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G48), .B2(new_n542), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n571), .B2(G86), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  AOI211_X1 g177(.A(KEYINPUT82), .B(new_n602), .C1(new_n568), .C2(new_n570), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n500), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  INV_X1    g182(.A(G47), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n515), .A2(new_n607), .B1(new_n608), .B2(new_n518), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT83), .Z(new_n613));
  XOR2_X1   g188(.A(KEYINPUT84), .B(KEYINPUT10), .Z(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT85), .B1(new_n571), .B2(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  AOI211_X1 g193(.A(new_n617), .B(new_n618), .C1(new_n568), .C2(new_n570), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n534), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G54), .B2(new_n542), .ZN(new_n624));
  OAI21_X1  g199(.A(G92), .B1(new_n578), .B2(new_n579), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n617), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n571), .A2(KEYINPUT85), .A3(G92), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(new_n614), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n620), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n613), .B1(G868), .B2(new_n629), .ZN(G284));
  OAI21_X1  g205(.A(new_n613), .B1(G868), .B2(new_n629), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  XNOR2_X1  g207(.A(G299), .B(KEYINPUT86), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT87), .ZN(G297));
  XNOR2_X1  g210(.A(new_n634), .B(KEYINPUT88), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n629), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g217(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT89), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT90), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT91), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n653));
  INV_X1    g228(.A(G123), .ZN(new_n654));
  INV_X1    g229(.A(G135), .ZN(new_n655));
  OAI221_X1 g230(.A(new_n653), .B1(new_n483), .B2(new_n654), .C1(new_n655), .C2(new_n486), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT92), .B(G2096), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n649), .A2(new_n651), .A3(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2435), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2438), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT93), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2443), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2446), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n670), .ZN(new_n672));
  XOR2_X1   g247(.A(G2451), .B(G2454), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT94), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n671), .B2(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(G14), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G401));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT96), .ZN(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2096), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n685), .B1(KEYINPUT97), .B2(KEYINPUT17), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n683), .A2(new_n684), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(KEYINPUT97), .C2(KEYINPUT17), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n686), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n699), .A2(new_n701), .A3(new_n703), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n706), .B(new_n707), .C1(new_n705), .C2(new_n704), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT98), .B(G1981), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n708), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT99), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n712), .B(new_n715), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  NOR2_X1   g292(.A1(G16), .A2(G24), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n610), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1986), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n481), .A2(new_n482), .A3(G119), .A4(G2105), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n482), .A3(G131), .A4(new_n462), .ZN(new_n724));
  OR2_X1    g299(.A1(G95), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(new_n721), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT100), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n720), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G23), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT33), .B(G1976), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G22), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G166), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1971), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G6), .ZN(new_n744));
  INV_X1    g319(.A(new_n599), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n571), .A2(G86), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT82), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n571), .A2(new_n600), .A3(G86), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(new_n743), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT32), .B(G1981), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT34), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT34), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n732), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT101), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(KEYINPUT36), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n732), .B1(new_n757), .B2(KEYINPUT36), .C1(new_n754), .C2(new_n755), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(new_n757), .B2(KEYINPUT36), .ZN(new_n761));
  OR2_X1    g336(.A1(G29), .A2(G33), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n481), .A2(new_n482), .A3(G139), .A4(new_n462), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G127), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n479), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2105), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n763), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT103), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT103), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n763), .A2(new_n767), .A3(new_n772), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n762), .B1(new_n774), .B2(new_n721), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT105), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n743), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n629), .B2(new_n743), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(G34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n464), .A2(new_n467), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2105), .ZN(new_n790));
  INV_X1    g365(.A(G137), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n470), .B1(new_n479), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(new_n462), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n788), .B1(new_n794), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT30), .B(G28), .Z(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(G29), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G2078), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT31), .B(G11), .Z(new_n803));
  NOR3_X1   g378(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G19), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n551), .B2(G16), .ZN(new_n806));
  AOI22_X1  g381(.A1(G1341), .A2(new_n806), .B1(new_n775), .B2(new_n776), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n795), .A2(new_n796), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT104), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n804), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n487), .A2(G29), .ZN(new_n811));
  INV_X1    g386(.A(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT106), .B1(new_n812), .B2(G29), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n812), .A2(KEYINPUT106), .A3(G29), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT29), .ZN(new_n816));
  INV_X1    g391(.A(G2090), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n811), .A2(new_n818), .A3(new_n813), .A4(new_n814), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT107), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n721), .A2(G26), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT28), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n481), .A2(new_n482), .A3(G128), .A4(G2105), .ZN(new_n824));
  OR2_X1    g399(.A1(G104), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n826));
  INV_X1    g401(.A(G140), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n826), .C1(new_n486), .C2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n828), .A2(new_n829), .A3(G29), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n828), .B2(G29), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n823), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G2067), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n820), .A2(new_n821), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n816), .A2(new_n819), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n837), .A2(KEYINPUT107), .A3(new_n817), .ZN(new_n838));
  OR2_X1    g413(.A1(G29), .A2(G32), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n481), .A2(new_n482), .A3(G141), .A4(new_n462), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n481), .A2(new_n482), .A3(G129), .A4(G2105), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n842));
  NAND3_X1  g417(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT26), .Z(new_n844));
  NAND4_X1  g419(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n839), .B1(new_n845), .B2(new_n721), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT27), .B(G1996), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n801), .A2(G2078), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n743), .A2(G5), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G171), .B2(new_n743), .ZN(new_n852));
  INV_X1    g427(.A(G1961), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(G1961), .B(new_n851), .C1(G171), .C2(new_n743), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n810), .A2(new_n836), .A3(new_n838), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n784), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n837), .A2(new_n817), .ZN(new_n859));
  NAND2_X1  g434(.A1(G299), .A2(G16), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n743), .A2(KEYINPUT23), .A3(G20), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT23), .ZN(new_n862));
  INV_X1    g437(.A(G20), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(G16), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G1956), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n859), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n858), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n743), .A2(G21), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(G168), .B2(new_n743), .ZN(new_n874));
  INV_X1    g449(.A(G1966), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n806), .A2(G1341), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n869), .A2(new_n870), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n872), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n721), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT109), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g457(.A(KEYINPUT108), .B(new_n859), .C1(new_n867), .C2(new_n868), .ZN(new_n883));
  INV_X1    g458(.A(new_n876), .ZN(new_n884));
  NOR4_X1   g459(.A1(new_n871), .A2(new_n883), .A3(new_n884), .A4(new_n877), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n886));
  INV_X1    g461(.A(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n761), .B1(new_n882), .B2(new_n888), .ZN(G311));
  INV_X1    g464(.A(new_n761), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n867), .A2(new_n868), .ZN(new_n892));
  INV_X1    g467(.A(new_n859), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT108), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n895), .A2(new_n878), .A3(new_n879), .A4(new_n858), .ZN(new_n896));
  NOR4_X1   g471(.A1(new_n896), .A2(KEYINPUT109), .A3(new_n881), .A4(new_n884), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n890), .B1(new_n891), .B2(new_n897), .ZN(G150));
  NAND2_X1  g473(.A1(new_n507), .A2(G67), .ZN(new_n899));
  NAND2_X1  g474(.A1(G80), .A2(G543), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n500), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G93), .ZN(new_n902));
  INV_X1    g477(.A(G55), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n515), .A2(new_n902), .B1(new_n903), .B2(new_n518), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(KEYINPUT111), .B(G860), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT112), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT37), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n620), .A2(new_n624), .A3(new_n628), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n637), .ZN(new_n916));
  XOR2_X1   g491(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n908), .B2(new_n909), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n905), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n918), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n914), .B1(new_n924), .B2(new_n911), .ZN(G145));
  INV_X1    g500(.A(KEYINPUT114), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n481), .A2(new_n482), .A3(G130), .A4(G2105), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n481), .A2(new_n482), .A3(G142), .A4(new_n462), .ZN(new_n928));
  OR2_X1    g503(.A1(G106), .A2(G2105), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n727), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n927), .A3(new_n928), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT113), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT113), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n644), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n644), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n932), .B2(new_n934), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n845), .B1(new_n771), .B2(new_n773), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT4), .B1(new_n463), .B2(G138), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n498), .B1(new_n946), .B2(G2105), .ZN(new_n947));
  INV_X1    g522(.A(new_n491), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n828), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n771), .A2(new_n773), .A3(new_n845), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n828), .B(G164), .ZN(new_n953));
  INV_X1    g528(.A(new_n951), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n944), .ZN(new_n955));
  AND4_X1   g530(.A1(new_n939), .A2(new_n943), .A3(new_n952), .A4(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n943), .A2(new_n939), .B1(new_n955), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n926), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n957), .A2(new_n926), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n656), .B(G160), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(G162), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n956), .B2(new_n957), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g542(.A(G868), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n749), .A2(G288), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n734), .A2(G305), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(G166), .ZN(new_n971));
  AOI21_X1  g546(.A(G166), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(G290), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G303), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n970), .A3(G166), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n610), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT42), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n639), .B(new_n923), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n616), .A2(new_n619), .A3(new_n615), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n614), .B1(new_n626), .B2(new_n627), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(new_n577), .A3(new_n585), .A4(new_n624), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n584), .B1(new_n583), .B2(new_n567), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT80), .B(new_n566), .C1(new_n581), .C2(new_n582), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n915), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n980), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT41), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n983), .A2(new_n624), .B1(new_n577), .B2(new_n585), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n915), .A2(new_n985), .A3(new_n986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n987), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n980), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n968), .B1(new_n979), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n979), .B2(new_n996), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n978), .B(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT115), .A3(new_n989), .A4(new_n995), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n968), .B1(new_n908), .B2(new_n909), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(KEYINPUT116), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(G295));
  INV_X1    g584(.A(new_n1005), .ZN(G331));
  AND2_X1   g585(.A1(new_n973), .A2(new_n977), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G301), .A2(G168), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G286), .A2(new_n541), .A3(new_n543), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n901), .A2(new_n904), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n551), .B1(new_n1016), .B2(new_n907), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n921), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n920), .A2(new_n922), .A3(new_n1013), .A4(new_n1012), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n993), .B2(new_n994), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n987), .B2(new_n984), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1011), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n987), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT41), .B1(new_n984), .B2(new_n987), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n988), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n978), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1029), .A3(new_n964), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1024), .A2(new_n1029), .A3(new_n1032), .A4(new_n964), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1034), .B(KEYINPUT44), .Z(G397));
  INV_X1    g610(.A(KEYINPUT126), .ZN(new_n1036));
  INV_X1    g611(.A(G1996), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n845), .B(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n828), .B(new_n833), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(G164), .B2(G1384), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G160), .A2(G40), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n933), .A2(new_n730), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n933), .A2(new_n730), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G290), .A2(G1986), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G290), .A2(G1986), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n790), .A2(new_n793), .A3(G40), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n493), .B1(new_n463), .B2(G126), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n497), .A2(new_n1063), .B1(new_n494), .B2(new_n462), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT45), .B(new_n1062), .C1(new_n1064), .C2(new_n491), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1042), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n875), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT50), .B1(new_n949), .B2(new_n1062), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(G1384), .C1(new_n947), .C2(new_n948), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n796), .B(new_n1061), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1071), .A3(G168), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1060), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1069), .B1(G164), .B2(G1384), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n949), .A2(KEYINPUT50), .A3(new_n1062), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1043), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1078), .A2(new_n796), .B1(new_n1066), .B2(new_n875), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT51), .B1(new_n1079), .B2(G168), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1059), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1066), .A2(new_n1084), .A3(G2078), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1061), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n853), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(new_n1066), .B2(G2078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1093));
  OAI211_X1 g668(.A(G8), .B(new_n1072), .C1(new_n1093), .C2(new_n1060), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1083), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n522), .A2(G8), .A3(new_n523), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT55), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n522), .A2(new_n1100), .A3(G8), .A4(new_n523), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1078), .A2(new_n817), .B1(new_n1066), .B2(new_n740), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1066), .A2(new_n740), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n817), .B(new_n1061), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(G8), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1981), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n599), .C1(new_n601), .C2(new_n603), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n515), .A2(new_n602), .ZN(new_n1113));
  OAI21_X1  g688(.A(G1981), .B1(new_n745), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G164), .A2(G1384), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1104), .B1(new_n1118), .B2(new_n1061), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1114), .A3(KEYINPUT49), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n593), .B1(new_n571), .B2(G87), .ZN(new_n1122));
  INV_X1    g697(.A(G87), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT81), .B(new_n1123), .C1(new_n568), .C2(new_n570), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT118), .A3(G1976), .A4(new_n592), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n590), .A2(G1976), .A3(new_n592), .A4(new_n594), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1119), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT52), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1126), .A2(new_n1133), .A3(new_n1119), .A4(new_n1129), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1121), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1110), .B(new_n1135), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1121), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1095), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1118), .A2(new_n1061), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1078), .A2(G1348), .B1(new_n1140), .B2(G2067), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n915), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n629), .A2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1086), .A2(new_n781), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n833), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n915), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1148), .B2(KEYINPUT60), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT56), .B(G2072), .Z(new_n1150));
  NOR2_X1   g725(.A1(new_n1066), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT120), .B(G1956), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1086), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n583), .B2(new_n567), .ZN(new_n1156));
  AOI211_X1 g731(.A(KEYINPUT121), .B(new_n566), .C1(new_n581), .C2(new_n582), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n576), .A2(KEYINPUT121), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n583), .A2(new_n1155), .A3(new_n567), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(KEYINPUT57), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT61), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT58), .B(G1341), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1145), .A2(new_n1164), .B1(new_n1066), .B2(G1996), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n551), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n551), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1153), .A2(new_n1158), .A3(new_n1171), .A4(new_n1161), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1149), .A2(new_n1163), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1153), .B1(new_n1161), .B2(new_n1158), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n629), .A2(new_n1141), .A3(KEYINPUT122), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT122), .B1(new_n629), .B2(new_n1141), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1177), .B2(new_n1162), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1139), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1085), .A2(new_n1087), .A3(G301), .A4(new_n1088), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1090), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT54), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1097), .A2(new_n1136), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1135), .A2(KEYINPUT119), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1109), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1121), .A2(new_n1131), .A3(new_n1186), .A4(new_n1134), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1121), .A2(new_n1132), .A3(new_n734), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1112), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1119), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1074), .A2(new_n1193), .A3(G286), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1184), .A2(new_n1138), .A3(new_n1187), .A4(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1137), .A2(new_n1138), .A3(G168), .A4(new_n1075), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1193), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1192), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1058), .B1(new_n1183), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1051), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1053), .A2(new_n1044), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1048), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1046), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n828), .A2(G2067), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1044), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(KEYINPUT124), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1210), .B(new_n1044), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n845), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1052), .B1(new_n1213), .B2(new_n1039), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1215), .B2(KEYINPUT46), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1044), .A2(new_n1037), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1215), .A2(KEYINPUT46), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1217), .B(new_n1218), .Z(new_n1219));
  NAND2_X1  g794(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT47), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1204), .A2(new_n1212), .A3(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1036), .B1(new_n1199), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1136), .A2(new_n1091), .A3(new_n1096), .A4(new_n1083), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1197), .A2(new_n1195), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1227), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1057), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1222), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1229), .A2(new_n1230), .A3(KEYINPUT126), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1223), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g807(.A(G401), .ZN(new_n1234));
  AND4_X1   g808(.A1(new_n460), .A2(new_n966), .A3(new_n694), .A4(new_n716), .ZN(new_n1235));
  AND4_X1   g809(.A1(KEYINPUT127), .A2(new_n1034), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(G401), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1237));
  AOI21_X1  g811(.A(KEYINPUT127), .B1(new_n1237), .B2(new_n1235), .ZN(new_n1238));
  NOR2_X1   g812(.A1(new_n1236), .A2(new_n1238), .ZN(G308));
  NAND3_X1  g813(.A1(new_n1034), .A2(new_n1235), .A3(new_n1234), .ZN(new_n1240));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g816(.A1(new_n1237), .A2(KEYINPUT127), .A3(new_n1235), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1242), .A2(new_n1243), .ZN(G225));
endmodule


