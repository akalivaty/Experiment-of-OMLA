

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751;

  AND2_X1 U373 ( .A1(n386), .A2(n385), .ZN(n384) );
  INV_X1 U374 ( .A(n702), .ZN(n351) );
  INV_X1 U375 ( .A(n626), .ZN(n350) );
  XNOR2_X1 U376 ( .A(n581), .B(KEYINPUT95), .ZN(n571) );
  XNOR2_X1 U377 ( .A(n579), .B(KEYINPUT109), .ZN(n541) );
  INV_X1 U378 ( .A(G128), .ZN(n412) );
  NAND2_X2 U379 ( .A1(n496), .A2(n479), .ZN(n497) );
  XNOR2_X2 U380 ( .A(n463), .B(n462), .ZN(n466) );
  NAND2_X1 U381 ( .A1(n351), .A2(n350), .ZN(n365) );
  BUF_X1 U382 ( .A(G953), .Z(n748) );
  XNOR2_X2 U383 ( .A(n740), .B(n416), .ZN(n485) );
  NOR2_X4 U384 ( .A1(n522), .A2(n574), .ZN(n659) );
  XNOR2_X1 U385 ( .A(n531), .B(n530), .ZN(n566) );
  OR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n358) );
  NAND2_X1 U387 ( .A1(n375), .A2(n356), .ZN(n564) );
  AND2_X1 U388 ( .A1(n566), .A2(n665), .ZN(n580) );
  BUF_X1 U389 ( .A(n566), .Z(n532) );
  XNOR2_X1 U390 ( .A(n402), .B(n401), .ZN(n669) );
  NOR2_X2 U391 ( .A1(G902), .A2(n714), .ZN(n439) );
  NOR2_X1 U392 ( .A1(n724), .A2(G902), .ZN(n402) );
  XNOR2_X1 U393 ( .A(n495), .B(n494), .ZN(n629) );
  BUF_X1 U394 ( .A(n599), .Z(n352) );
  BUF_X1 U395 ( .A(n680), .Z(n353) );
  XNOR2_X1 U396 ( .A(n570), .B(n569), .ZN(n680) );
  AND2_X1 U397 ( .A1(n386), .A2(KEYINPUT85), .ZN(n354) );
  BUF_X1 U398 ( .A(n351), .Z(n355) );
  BUF_X1 U399 ( .A(n713), .Z(n723) );
  XNOR2_X1 U400 ( .A(G113), .B(G101), .ZN(n471) );
  XNOR2_X1 U401 ( .A(G119), .B(G116), .ZN(n470) );
  NAND2_X1 U402 ( .A1(n366), .A2(KEYINPUT2), .ZN(n386) );
  XNOR2_X1 U403 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  XOR2_X1 U404 ( .A(G137), .B(G140), .Z(n406) );
  XNOR2_X1 U405 ( .A(n379), .B(G146), .ZN(n464) );
  INV_X1 U406 ( .A(G125), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n371), .B(n505), .ZN(n602) );
  NAND2_X1 U408 ( .A1(n504), .A2(n503), .ZN(n371) );
  INV_X1 U409 ( .A(n592), .ZN(n378) );
  XNOR2_X1 U410 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U411 ( .A1(n713), .A2(G210), .ZN(n367) );
  XNOR2_X1 U412 ( .A(n640), .B(n642), .ZN(n643) );
  AND2_X1 U413 ( .A1(n633), .A2(n632), .ZN(n728) );
  INV_X1 U414 ( .A(G237), .ZN(n478) );
  XNOR2_X1 U415 ( .A(KEYINPUT71), .B(KEYINPUT93), .ZN(n469) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n426) );
  INV_X1 U417 ( .A(n626), .ZN(n385) );
  XOR2_X1 U418 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n462) );
  NAND2_X1 U419 ( .A1(n602), .A2(n509), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n430), .B(n396), .ZN(n741) );
  XNOR2_X1 U421 ( .A(G134), .B(G116), .ZN(n441) );
  INV_X1 U422 ( .A(G146), .ZN(n416) );
  XNOR2_X1 U423 ( .A(G110), .B(G107), .ZN(n407) );
  BUF_X1 U424 ( .A(n537), .Z(n581) );
  XNOR2_X1 U425 ( .A(G143), .B(G113), .ZN(n423) );
  XNOR2_X1 U426 ( .A(n560), .B(n559), .ZN(n599) );
  NAND2_X1 U427 ( .A1(n378), .A2(n377), .ZN(n375) );
  NOR2_X1 U428 ( .A1(n539), .A2(KEYINPUT66), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n367), .B(n643), .ZN(n644) );
  XNOR2_X1 U430 ( .A(n712), .B(n363), .ZN(G75) );
  INV_X1 U431 ( .A(KEYINPUT53), .ZN(n363) );
  AND2_X1 U432 ( .A1(n372), .A2(n361), .ZN(n356) );
  NOR2_X1 U433 ( .A1(n575), .A2(n514), .ZN(n357) );
  XOR2_X1 U434 ( .A(KEYINPUT65), .B(KEYINPUT4), .Z(n359) );
  XOR2_X1 U435 ( .A(KEYINPUT84), .B(n700), .Z(n360) );
  AND2_X1 U436 ( .A1(n376), .A2(n588), .ZN(n361) );
  OR2_X1 U437 ( .A1(n625), .A2(KEYINPUT2), .ZN(n362) );
  NOR2_X1 U438 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U439 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U440 ( .A(n485), .B(n417), .ZN(n647) );
  INV_X1 U441 ( .A(n629), .ZN(n496) );
  NAND2_X1 U442 ( .A1(n384), .A2(n362), .ZN(n368) );
  XNOR2_X2 U443 ( .A(n364), .B(n521), .ZN(n558) );
  NAND2_X1 U444 ( .A1(n519), .A2(n520), .ZN(n364) );
  XNOR2_X1 U445 ( .A(n467), .B(n468), .ZN(n477) );
  NOR2_X2 U446 ( .A1(n680), .A2(n571), .ZN(n573) );
  NAND2_X1 U447 ( .A1(n354), .A2(n365), .ZN(n369) );
  INV_X1 U448 ( .A(n701), .ZN(n366) );
  XNOR2_X1 U449 ( .A(n580), .B(KEYINPUT110), .ZN(n568) );
  NAND2_X2 U450 ( .A1(n369), .A2(n368), .ZN(n713) );
  XNOR2_X1 U451 ( .A(n381), .B(n565), .ZN(n380) );
  XNOR2_X2 U452 ( .A(n370), .B(n511), .ZN(n537) );
  NAND2_X1 U453 ( .A1(n638), .A2(n564), .ZN(n381) );
  NAND2_X1 U454 ( .A1(n592), .A2(KEYINPUT66), .ZN(n372) );
  XNOR2_X2 U455 ( .A(n373), .B(KEYINPUT32), .ZN(n638) );
  OR2_X2 U456 ( .A1(n592), .A2(n374), .ZN(n373) );
  NAND2_X1 U457 ( .A1(n563), .A2(n562), .ZN(n374) );
  XNOR2_X2 U458 ( .A(n538), .B(KEYINPUT22), .ZN(n592) );
  NAND2_X1 U459 ( .A1(n539), .A2(KEYINPUT66), .ZN(n376) );
  NOR2_X2 U460 ( .A1(n639), .A2(n380), .ZN(n578) );
  XNOR2_X2 U461 ( .A(n382), .B(KEYINPUT35), .ZN(n639) );
  NAND2_X1 U462 ( .A1(n383), .A2(n577), .ZN(n382) );
  XNOR2_X1 U463 ( .A(n573), .B(n572), .ZN(n383) );
  XNOR2_X2 U464 ( .A(n467), .B(n415), .ZN(n740) );
  XNOR2_X2 U465 ( .A(n440), .B(n359), .ZN(n467) );
  XNOR2_X2 U466 ( .A(n413), .B(n412), .ZN(n440) );
  NOR2_X1 U467 ( .A1(n571), .A2(n513), .ZN(n583) );
  INV_X1 U468 ( .A(KEYINPUT107), .ZN(n586) );
  XNOR2_X1 U469 ( .A(n587), .B(n586), .ZN(n593) );
  BUF_X1 U470 ( .A(n461), .Z(n633) );
  XOR2_X1 U471 ( .A(KEYINPUT98), .B(G110), .Z(n388) );
  XNOR2_X1 U472 ( .A(G128), .B(G119), .ZN(n387) );
  XNOR2_X1 U473 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n390) );
  XNOR2_X1 U475 ( .A(KEYINPUT76), .B(KEYINPUT24), .ZN(n389) );
  XNOR2_X1 U476 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U477 ( .A(n392), .B(n391), .Z(n395) );
  XNOR2_X2 U478 ( .A(KEYINPUT64), .B(G953), .ZN(n461) );
  INV_X1 U479 ( .A(n461), .ZN(n743) );
  NAND2_X1 U480 ( .A1(n743), .A2(G234), .ZN(n393) );
  XOR2_X1 U481 ( .A(KEYINPUT8), .B(n393), .Z(n447) );
  NAND2_X1 U482 ( .A1(G221), .A2(n447), .ZN(n394) );
  XNOR2_X1 U483 ( .A(n394), .B(n395), .ZN(n397) );
  XOR2_X1 U484 ( .A(n464), .B(KEYINPUT10), .Z(n430) );
  INV_X1 U485 ( .A(n406), .ZN(n396) );
  XNOR2_X1 U486 ( .A(n397), .B(n741), .ZN(n724) );
  NAND2_X1 U487 ( .A1(n626), .A2(G234), .ZN(n398) );
  XNOR2_X1 U488 ( .A(n398), .B(KEYINPUT20), .ZN(n403) );
  NAND2_X1 U489 ( .A1(n403), .A2(G217), .ZN(n400) );
  XOR2_X1 U490 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n399) );
  XNOR2_X1 U491 ( .A(n400), .B(n399), .ZN(n401) );
  NAND2_X1 U492 ( .A1(G221), .A2(n403), .ZN(n404) );
  XOR2_X1 U493 ( .A(KEYINPUT21), .B(n404), .Z(n668) );
  XNOR2_X1 U494 ( .A(n668), .B(KEYINPUT99), .ZN(n535) );
  INV_X1 U495 ( .A(n535), .ZN(n405) );
  AND2_X1 U496 ( .A1(n669), .A2(n405), .ZN(n665) );
  INV_X1 U497 ( .A(n665), .ZN(n422) );
  XOR2_X1 U498 ( .A(KEYINPUT96), .B(n406), .Z(n408) );
  XNOR2_X1 U499 ( .A(n407), .B(G104), .ZN(n475) );
  XNOR2_X1 U500 ( .A(n408), .B(n475), .ZN(n411) );
  INV_X1 U501 ( .A(G227), .ZN(n745) );
  OR2_X1 U502 ( .A1(n633), .A2(n745), .ZN(n409) );
  XNOR2_X1 U503 ( .A(n409), .B(G101), .ZN(n410) );
  XNOR2_X1 U504 ( .A(n411), .B(n410), .ZN(n417) );
  XNOR2_X2 U505 ( .A(G143), .B(KEYINPUT81), .ZN(n413) );
  INV_X1 U506 ( .A(KEYINPUT69), .ZN(n414) );
  XNOR2_X1 U507 ( .A(n414), .B(G131), .ZN(n431) );
  XNOR2_X1 U508 ( .A(n431), .B(G134), .ZN(n415) );
  OR2_X2 U509 ( .A1(n647), .A2(G902), .ZN(n420) );
  INV_X1 U510 ( .A(KEYINPUT70), .ZN(n418) );
  XNOR2_X1 U511 ( .A(n418), .B(G469), .ZN(n419) );
  XNOR2_X2 U512 ( .A(n420), .B(n419), .ZN(n531) );
  BUF_X1 U513 ( .A(n531), .Z(n421) );
  NOR2_X2 U514 ( .A1(n422), .A2(n421), .ZN(n512) );
  XNOR2_X1 U515 ( .A(n512), .B(KEYINPUT111), .ZN(n518) );
  INV_X1 U516 ( .A(n518), .ZN(n484) );
  XOR2_X1 U517 ( .A(G140), .B(G104), .Z(n424) );
  XOR2_X1 U518 ( .A(n424), .B(n423), .Z(n435) );
  XNOR2_X2 U519 ( .A(KEYINPUT73), .B(n358), .ZN(n486) );
  NAND2_X1 U520 ( .A1(G214), .A2(n486), .ZN(n428) );
  XNOR2_X1 U521 ( .A(G122), .B(KEYINPUT102), .ZN(n425) );
  XNOR2_X1 U522 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U524 ( .A(n429), .B(KEYINPUT11), .Z(n433) );
  XNOR2_X1 U525 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U526 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U527 ( .A(n435), .B(n434), .ZN(n714) );
  XNOR2_X1 U528 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n437) );
  INV_X1 U529 ( .A(G475), .ZN(n436) );
  XNOR2_X2 U530 ( .A(n439), .B(n438), .ZN(n575) );
  INV_X1 U531 ( .A(n575), .ZN(n522) );
  XNOR2_X1 U532 ( .A(n441), .B(KEYINPUT7), .ZN(n445) );
  XOR2_X1 U533 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n443) );
  XNOR2_X1 U534 ( .A(G107), .B(G122), .ZN(n442) );
  XNOR2_X1 U535 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U536 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U537 ( .A(n440), .B(n446), .ZN(n449) );
  NAND2_X1 U538 ( .A1(G217), .A2(n447), .ZN(n448) );
  XNOR2_X1 U539 ( .A(n449), .B(n448), .ZN(n719) );
  INV_X1 U540 ( .A(G902), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n719), .A2(n479), .ZN(n451) );
  INV_X1 U542 ( .A(G478), .ZN(n450) );
  XNOR2_X2 U543 ( .A(n451), .B(n450), .ZN(n574) );
  NAND2_X1 U544 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U545 ( .A(n452), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U546 ( .A1(G952), .A2(n455), .ZN(n453) );
  XNOR2_X1 U547 ( .A(KEYINPUT94), .B(n453), .ZN(n698) );
  INV_X1 U548 ( .A(n698), .ZN(n454) );
  INV_X1 U549 ( .A(n748), .ZN(n729) );
  NAND2_X1 U550 ( .A1(n454), .A2(n729), .ZN(n508) );
  AND2_X1 U551 ( .A1(G902), .A2(n455), .ZN(n506) );
  NAND2_X1 U552 ( .A1(n633), .A2(n506), .ZN(n456) );
  OR2_X1 U553 ( .A1(G900), .A2(n456), .ZN(n457) );
  NAND2_X1 U554 ( .A1(n508), .A2(n457), .ZN(n523) );
  INV_X1 U555 ( .A(n523), .ZN(n458) );
  NOR2_X1 U556 ( .A1(n574), .A2(n458), .ZN(n459) );
  NAND2_X1 U557 ( .A1(n522), .A2(n459), .ZN(n482) );
  INV_X1 U558 ( .A(G224), .ZN(n460) );
  OR2_X2 U559 ( .A1(n461), .A2(n460), .ZN(n463) );
  XNOR2_X1 U560 ( .A(n464), .B(KEYINPUT77), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n470), .B(n469), .ZN(n473) );
  XNOR2_X1 U563 ( .A(n471), .B(KEYINPUT3), .ZN(n472) );
  XNOR2_X1 U564 ( .A(n473), .B(n472), .ZN(n492) );
  XNOR2_X1 U565 ( .A(KEYINPUT16), .B(G122), .ZN(n474) );
  XNOR2_X1 U566 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U567 ( .A(n492), .B(n476), .ZN(n734) );
  XNOR2_X1 U568 ( .A(n477), .B(n734), .ZN(n640) );
  NAND2_X1 U569 ( .A1(n640), .A2(n626), .ZN(n481) );
  NAND2_X1 U570 ( .A1(n479), .A2(n478), .ZN(n498) );
  NAND2_X1 U571 ( .A1(n498), .A2(G210), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n481), .B(n480), .ZN(n502) );
  BUF_X1 U573 ( .A(n502), .Z(n551) );
  NOR2_X1 U574 ( .A1(n482), .A2(n551), .ZN(n483) );
  NAND2_X1 U575 ( .A1(n484), .A2(n483), .ZN(n501) );
  INV_X1 U576 ( .A(n485), .ZN(n495) );
  XOR2_X1 U577 ( .A(KEYINPUT5), .B(G137), .Z(n488) );
  NAND2_X1 U578 ( .A1(n486), .A2(G210), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n488), .B(n487), .ZN(n491) );
  XNOR2_X1 U580 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U581 ( .A(n489), .B(KEYINPUT72), .ZN(n490) );
  XNOR2_X1 U582 ( .A(n491), .B(n490), .ZN(n493) );
  XNOR2_X1 U583 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X2 U584 ( .A(n497), .B(G472), .ZN(n579) );
  AND2_X1 U585 ( .A1(n498), .A2(G214), .ZN(n681) );
  NOR2_X1 U586 ( .A1(n541), .A2(n681), .ZN(n499) );
  XNOR2_X1 U587 ( .A(n499), .B(KEYINPUT30), .ZN(n519) );
  INV_X1 U588 ( .A(n519), .ZN(n500) );
  NOR2_X1 U589 ( .A1(n501), .A2(n500), .ZN(n612) );
  XOR2_X1 U590 ( .A(G143), .B(n612), .Z(G45) );
  INV_X1 U591 ( .A(n502), .ZN(n504) );
  INV_X1 U592 ( .A(n681), .ZN(n503) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n505) );
  NOR2_X1 U594 ( .A1(G898), .A2(n729), .ZN(n735) );
  NAND2_X1 U595 ( .A1(n506), .A2(n735), .ZN(n507) );
  NAND2_X1 U596 ( .A1(n508), .A2(n507), .ZN(n509) );
  INV_X1 U597 ( .A(KEYINPUT68), .ZN(n510) );
  XNOR2_X1 U598 ( .A(n510), .B(KEYINPUT0), .ZN(n511) );
  INV_X1 U599 ( .A(n579), .ZN(n671) );
  NAND2_X1 U600 ( .A1(n512), .A2(n671), .ZN(n513) );
  INV_X1 U601 ( .A(n574), .ZN(n514) );
  NAND2_X1 U602 ( .A1(n583), .A2(n357), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n515), .B(G104), .ZN(G6) );
  INV_X1 U604 ( .A(KEYINPUT38), .ZN(n516) );
  XNOR2_X1 U605 ( .A(n551), .B(n516), .ZN(n546) );
  INV_X1 U606 ( .A(n546), .ZN(n682) );
  NAND2_X1 U607 ( .A1(n682), .A2(n523), .ZN(n517) );
  NOR2_X1 U608 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U609 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n521) );
  XNOR2_X1 U610 ( .A(n659), .B(KEYINPUT106), .ZN(n584) );
  NAND2_X1 U611 ( .A1(n558), .A2(n584), .ZN(n622) );
  XNOR2_X1 U612 ( .A(n622), .B(G134), .ZN(G36) );
  NAND2_X1 U613 ( .A1(n668), .A2(n523), .ZN(n524) );
  OR2_X1 U614 ( .A1(n669), .A2(n524), .ZN(n540) );
  NOR2_X1 U615 ( .A1(n540), .A2(n681), .ZN(n525) );
  NAND2_X1 U616 ( .A1(n525), .A2(n357), .ZN(n526) );
  XNOR2_X2 U617 ( .A(n579), .B(KEYINPUT6), .ZN(n589) );
  NOR2_X1 U618 ( .A1(n526), .A2(n589), .ZN(n549) );
  INV_X1 U619 ( .A(n551), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n549), .A2(n527), .ZN(n529) );
  XOR2_X1 U621 ( .A(KEYINPUT90), .B(KEYINPUT36), .Z(n528) );
  XNOR2_X1 U622 ( .A(n529), .B(n528), .ZN(n533) );
  XNOR2_X1 U623 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n530) );
  NAND2_X1 U624 ( .A1(n533), .A2(n532), .ZN(n614) );
  XOR2_X1 U625 ( .A(G125), .B(KEYINPUT37), .Z(n534) );
  XNOR2_X1 U626 ( .A(n614), .B(n534), .ZN(G27) );
  NAND2_X1 U627 ( .A1(n575), .A2(n574), .ZN(n684) );
  NOR2_X1 U628 ( .A1(n684), .A2(n535), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U630 ( .A(n532), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n561), .A2(n541), .ZN(n539) );
  INV_X1 U632 ( .A(n669), .ZN(n588) );
  XNOR2_X1 U633 ( .A(n564), .B(G110), .ZN(G12) );
  NOR2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n542), .B(KEYINPUT28), .ZN(n544) );
  XOR2_X1 U636 ( .A(KEYINPUT112), .B(n421), .Z(n543) );
  NAND2_X1 U637 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U638 ( .A(n545), .B(KEYINPUT113), .ZN(n603) );
  OR2_X1 U639 ( .A1(n546), .A2(n681), .ZN(n686) );
  OR2_X1 U640 ( .A1(n684), .A2(n686), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT41), .ZN(n678) );
  NAND2_X1 U642 ( .A1(n603), .A2(n678), .ZN(n548) );
  XNOR2_X1 U643 ( .A(n548), .B(KEYINPUT42), .ZN(n598) );
  XNOR2_X1 U644 ( .A(n598), .B(G137), .ZN(G39) );
  NAND2_X1 U645 ( .A1(n549), .A2(n561), .ZN(n550) );
  XNOR2_X1 U646 ( .A(n550), .B(KEYINPUT43), .ZN(n552) );
  NAND2_X1 U647 ( .A1(n552), .A2(n551), .ZN(n621) );
  XNOR2_X1 U648 ( .A(n621), .B(G140), .ZN(G42) );
  NAND2_X1 U649 ( .A1(n583), .A2(n659), .ZN(n557) );
  XOR2_X1 U650 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n554) );
  XNOR2_X1 U651 ( .A(G107), .B(KEYINPUT26), .ZN(n553) );
  XNOR2_X1 U652 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U653 ( .A(KEYINPUT116), .B(n555), .Z(n556) );
  XNOR2_X1 U654 ( .A(n557), .B(n556), .ZN(G9) );
  NAND2_X1 U655 ( .A1(n558), .A2(n357), .ZN(n560) );
  XNOR2_X1 U656 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n559) );
  XNOR2_X1 U657 ( .A(n352), .B(G131), .ZN(G33) );
  INV_X1 U658 ( .A(KEYINPUT89), .ZN(n565) );
  NOR2_X1 U659 ( .A1(n561), .A2(n669), .ZN(n563) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT80), .ZN(n562) );
  INV_X1 U661 ( .A(n589), .ZN(n567) );
  NAND2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U663 ( .A(KEYINPUT33), .ZN(n569) );
  XOR2_X1 U664 ( .A(KEYINPUT79), .B(KEYINPUT34), .Z(n572) );
  NOR2_X1 U665 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U666 ( .A(n576), .B(KEYINPUT78), .ZN(n577) );
  XNOR2_X1 U667 ( .A(n578), .B(KEYINPUT44), .ZN(n596) );
  AND2_X1 U668 ( .A1(n579), .A2(n580), .ZN(n675) );
  NAND2_X1 U669 ( .A1(n675), .A2(n581), .ZN(n582) );
  XNOR2_X1 U670 ( .A(n582), .B(KEYINPUT31), .ZN(n660) );
  NOR2_X1 U671 ( .A1(n660), .A2(n583), .ZN(n585) );
  NOR2_X2 U672 ( .A1(n584), .A2(n357), .ZN(n687) );
  XOR2_X1 U673 ( .A(KEYINPUT83), .B(n687), .Z(n604) );
  NOR2_X1 U674 ( .A1(n585), .A2(n604), .ZN(n587) );
  NOR2_X1 U675 ( .A1(n532), .A2(n588), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n652) );
  NOR2_X1 U678 ( .A1(n593), .A2(n652), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n594), .B(KEYINPUT108), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X2 U681 ( .A(n597), .B(KEYINPUT45), .ZN(n699) );
  NAND2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n601) );
  XNOR2_X1 U683 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n600) );
  XNOR2_X1 U684 ( .A(n601), .B(n600), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n653) );
  NOR2_X1 U686 ( .A1(n604), .A2(n653), .ZN(n607) );
  INV_X1 U687 ( .A(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n605), .A2(KEYINPUT82), .ZN(n606) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n687), .A2(KEYINPUT82), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n608), .A2(KEYINPUT47), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n653), .A2(n609), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n687), .A2(KEYINPUT82), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT48), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X2 U701 ( .A1(n624), .A2(n623), .ZN(n742) );
  NAND2_X2 U702 ( .A1(n699), .A2(n742), .ZN(n701) );
  NOR2_X1 U703 ( .A1(n701), .A2(KEYINPUT85), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n713), .A2(G472), .ZN(n631) );
  XNOR2_X1 U705 ( .A(KEYINPUT92), .B(KEYINPUT62), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n634) );
  INV_X1 U708 ( .A(G952), .ZN(n632) );
  NOR2_X2 U709 ( .A1(n634), .A2(n728), .ZN(n636) );
  XNOR2_X1 U710 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n636), .B(n635), .ZN(G57) );
  XOR2_X1 U712 ( .A(G119), .B(KEYINPUT127), .Z(n637) );
  XNOR2_X1 U713 ( .A(n638), .B(n637), .ZN(G21) );
  XOR2_X1 U714 ( .A(n639), .B(G122), .Z(G24) );
  XNOR2_X1 U715 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n641) );
  XOR2_X1 U716 ( .A(n641), .B(KEYINPUT55), .Z(n642) );
  NOR2_X2 U717 ( .A1(n644), .A2(n728), .ZN(n646) );
  XNOR2_X1 U718 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n646), .B(n645), .ZN(G51) );
  NAND2_X1 U720 ( .A1(n723), .A2(G469), .ZN(n650) );
  XOR2_X1 U721 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n648) );
  XNOR2_X1 U722 ( .A(n647), .B(n648), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U724 ( .A1(n651), .A2(n728), .ZN(G54) );
  XOR2_X1 U725 ( .A(G101), .B(n652), .Z(G3) );
  XOR2_X1 U726 ( .A(G128), .B(KEYINPUT29), .Z(n655) );
  INV_X1 U727 ( .A(n653), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n656), .A2(n659), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(G30) );
  NAND2_X1 U730 ( .A1(n656), .A2(n357), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(G146), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n660), .A2(n357), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(G113), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(KEYINPUT118), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G116), .B(n662), .ZN(G18) );
  INV_X1 U737 ( .A(n678), .ZN(n663) );
  NOR2_X1 U738 ( .A1(n353), .A2(n663), .ZN(n664) );
  NOR2_X1 U739 ( .A1(n664), .A2(n748), .ZN(n711) );
  NOR2_X1 U740 ( .A1(n532), .A2(n665), .ZN(n667) );
  XOR2_X1 U741 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U744 ( .A(KEYINPUT49), .B(n670), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U748 ( .A(KEYINPUT51), .B(n677), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n694) );
  INV_X1 U750 ( .A(n353), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n682), .A2(n503), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT120), .B(n685), .Z(n690) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(KEYINPUT121), .B(n688), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U759 ( .A(n695), .B(KEYINPUT122), .Z(n696) );
  XNOR2_X1 U760 ( .A(KEYINPUT52), .B(n696), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n709) );
  BUF_X1 U762 ( .A(n699), .Z(n700) );
  NOR2_X1 U763 ( .A1(n360), .A2(KEYINPUT2), .ZN(n705) );
  BUF_X1 U764 ( .A(n701), .Z(n702) );
  NAND2_X1 U765 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n355), .A2(n703), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n742), .A2(KEYINPUT2), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U770 ( .A1(n713), .A2(G475), .ZN(n716) );
  XOR2_X1 U771 ( .A(n714), .B(KEYINPUT59), .Z(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X2 U773 ( .A1(n717), .A2(n728), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U775 ( .A1(n723), .A2(G478), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n719), .B(KEYINPUT123), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n728), .A2(n722), .ZN(G63) );
  NAND2_X1 U779 ( .A1(n723), .A2(G217), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n724), .B(KEYINPUT124), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U783 ( .A1(n700), .A2(n729), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n748), .A2(G224), .ZN(n730) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n731), .A2(G898), .ZN(n732) );
  NAND2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n738) );
  XOR2_X1 U788 ( .A(KEYINPUT125), .B(n734), .Z(n736) );
  NOR2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U791 ( .A(KEYINPUT126), .B(n739), .ZN(G69) );
  XNOR2_X1 U792 ( .A(n740), .B(n741), .ZN(n746) );
  XNOR2_X1 U793 ( .A(n742), .B(n746), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n751) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n747), .A2(G900), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n751), .A2(n750), .ZN(G72) );
endmodule

