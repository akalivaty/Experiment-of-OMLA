

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  XNOR2_X1 U322 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U323 ( .A(n314), .B(n290), .ZN(n300) );
  XNOR2_X1 U324 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n468) );
  XNOR2_X1 U325 ( .A(n329), .B(n328), .ZN(n332) );
  XNOR2_X1 U326 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n380) );
  XNOR2_X1 U327 ( .A(n484), .B(KEYINPUT97), .ZN(n492) );
  XNOR2_X1 U328 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U329 ( .A(n307), .B(n306), .Z(n576) );
  AND2_X1 U330 ( .A1(G229GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U331 ( .A(n422), .B(n365), .Z(n291) );
  XNOR2_X1 U332 ( .A(n364), .B(n327), .ZN(n328) );
  XNOR2_X1 U333 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n368) );
  INV_X1 U334 ( .A(G197GAT), .ZN(n386) );
  INV_X1 U335 ( .A(KEYINPUT67), .ZN(n353) );
  XNOR2_X1 U336 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U337 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U338 ( .A(n531), .B(n468), .ZN(n478) );
  XNOR2_X1 U339 ( .A(n389), .B(n388), .ZN(n429) );
  XNOR2_X1 U340 ( .A(n393), .B(n355), .ZN(n359) );
  XNOR2_X1 U341 ( .A(n341), .B(n340), .ZN(n345) );
  INV_X1 U342 ( .A(n492), .ZN(n493) );
  INV_X1 U343 ( .A(KEYINPUT120), .ZN(n457) );
  XNOR2_X1 U344 ( .A(n346), .B(KEYINPUT65), .ZN(n347) );
  NOR2_X1 U345 ( .A1(n418), .A2(n529), .ZN(n575) );
  XNOR2_X1 U346 ( .A(n458), .B(n457), .ZN(n571) );
  XNOR2_X1 U347 ( .A(n370), .B(n347), .ZN(n560) );
  XNOR2_X1 U348 ( .A(n366), .B(n291), .ZN(n568) );
  XNOR2_X1 U349 ( .A(n372), .B(n371), .ZN(n553) );
  XNOR2_X1 U350 ( .A(n465), .B(G190GAT), .ZN(n466) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U352 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(G1GAT), .B(G113GAT), .Z(n293) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G197GAT), .ZN(n292) );
  XNOR2_X1 U355 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U356 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n295) );
  XNOR2_X1 U357 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n294) );
  XNOR2_X1 U358 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n297), .B(n296), .ZN(n307) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U362 ( .A(n299), .B(n298), .ZN(n301) );
  XOR2_X1 U363 ( .A(G22GAT), .B(G15GAT), .Z(n314) );
  XOR2_X1 U364 ( .A(n302), .B(KEYINPUT29), .Z(n305) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n303), .B(KEYINPUT7), .ZN(n361) );
  XNOR2_X1 U367 ( .A(n361), .B(KEYINPUT30), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U369 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n398) );
  XOR2_X1 U370 ( .A(KEYINPUT78), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n382) );
  XOR2_X1 U373 ( .A(G1GAT), .B(G127GAT), .Z(n405) );
  XOR2_X1 U374 ( .A(n382), .B(n405), .Z(n316) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U376 ( .A(n310), .B(KEYINPUT13), .ZN(n335) );
  XOR2_X1 U377 ( .A(G57GAT), .B(n335), .Z(n312) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U379 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U381 ( .A(n316), .B(n315), .ZN(n324) );
  XOR2_X1 U382 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n318) );
  XNOR2_X1 U383 ( .A(G155GAT), .B(KEYINPUT12), .ZN(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U385 ( .A(G64GAT), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U386 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U388 ( .A(n322), .B(n321), .Z(n323) );
  XOR2_X1 U389 ( .A(n324), .B(n323), .Z(n565) );
  XOR2_X1 U390 ( .A(KEYINPUT111), .B(n565), .Z(n570) );
  XOR2_X1 U391 ( .A(G92GAT), .B(KEYINPUT72), .Z(n326) );
  XNOR2_X1 U392 ( .A(G204GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U393 ( .A(n326), .B(n325), .ZN(n329) );
  XNOR2_X1 U394 ( .A(G99GAT), .B(G106GAT), .ZN(n364) );
  NAND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  INV_X1 U396 ( .A(n332), .ZN(n330) );
  NAND2_X1 U397 ( .A1(n330), .A2(KEYINPUT31), .ZN(n334) );
  INV_X1 U398 ( .A(KEYINPUT31), .ZN(n331) );
  NAND2_X1 U399 ( .A1(n332), .A2(n331), .ZN(n333) );
  NAND2_X1 U400 ( .A1(n334), .A2(n333), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n335), .B(KEYINPUT75), .ZN(n339) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(KEYINPUT71), .Z(n337) );
  XNOR2_X1 U403 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n336) );
  XOR2_X1 U404 ( .A(n337), .B(n336), .Z(n338) );
  XNOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n342), .B(KEYINPUT73), .ZN(n383) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(G148GAT), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n343), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U409 ( .A(n383), .B(n399), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n370) );
  INV_X1 U411 ( .A(KEYINPUT41), .ZN(n346) );
  INV_X1 U412 ( .A(n576), .ZN(n558) );
  AND2_X1 U413 ( .A1(n560), .A2(n558), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n348), .B(KEYINPUT46), .ZN(n349) );
  NOR2_X1 U415 ( .A1(n570), .A2(n349), .ZN(n350) );
  XNOR2_X1 U416 ( .A(KEYINPUT112), .B(n350), .ZN(n367) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G218GAT), .Z(n352) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n393) );
  NAND2_X1 U420 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XOR2_X1 U421 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n357) );
  XNOR2_X1 U422 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n363) );
  XNOR2_X1 U425 ( .A(G29GAT), .B(G134GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n360), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U427 ( .A(n361), .B(n409), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n366) );
  XOR2_X1 U429 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  INV_X1 U430 ( .A(n364), .ZN(n365) );
  INV_X1 U431 ( .A(n568), .ZN(n371) );
  NAND2_X1 U432 ( .A1(n367), .A2(n371), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n379) );
  INV_X1 U434 ( .A(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT36), .B(n553), .ZN(n587) );
  INV_X1 U436 ( .A(n565), .ZN(n584) );
  NOR2_X1 U437 ( .A1(n587), .A2(n584), .ZN(n374) );
  XNOR2_X1 U438 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  NAND2_X1 U440 ( .A1(n370), .A2(n375), .ZN(n376) );
  NOR2_X1 U441 ( .A1(n558), .A2(n376), .ZN(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT115), .B(n377), .ZN(n378) );
  AND2_X1 U443 ( .A1(n379), .A2(n378), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n539) );
  XOR2_X1 U445 ( .A(n383), .B(n382), .Z(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n385) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n448) );
  XNOR2_X1 U449 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n387) );
  XOR2_X1 U450 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n388) );
  XNOR2_X1 U451 ( .A(n448), .B(n429), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U453 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XOR2_X1 U455 ( .A(n395), .B(n394), .Z(n531) );
  INV_X1 U456 ( .A(n531), .ZN(n396) );
  NOR2_X1 U457 ( .A1(n539), .A2(n396), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n418) );
  XOR2_X1 U459 ( .A(G113GAT), .B(KEYINPUT0), .Z(n449) );
  XOR2_X1 U460 ( .A(n399), .B(n449), .Z(n401) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U464 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U466 ( .A(n404), .B(KEYINPUT92), .Z(n407) );
  XNOR2_X1 U467 ( .A(G162GAT), .B(n405), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U469 ( .A(n408), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U470 ( .A(n409), .B(KEYINPUT91), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U473 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U476 ( .A(G141GAT), .B(n416), .Z(n433) );
  XOR2_X1 U477 ( .A(n417), .B(n433), .Z(n475) );
  XNOR2_X1 U478 ( .A(KEYINPUT93), .B(n475), .ZN(n529) );
  XOR2_X1 U479 ( .A(G148GAT), .B(G211GAT), .Z(n420) );
  XNOR2_X1 U480 ( .A(G218GAT), .B(G106GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n421), .B(G78GAT), .Z(n424) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n426) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n428), .B(n427), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(KEYINPUT22), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n479) );
  NAND2_X1 U492 ( .A1(n575), .A2(n479), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n434), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U494 ( .A(G120GAT), .B(G176GAT), .Z(n436) );
  XNOR2_X1 U495 ( .A(G134GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n438) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(G127GAT), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n445) );
  XOR2_X1 U501 ( .A(G71GAT), .B(G183GAT), .Z(n442) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(KEYINPUT20), .B(n443), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT66), .B(KEYINPUT85), .Z(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n453) );
  XOR2_X1 U509 ( .A(n449), .B(n448), .Z(n451) );
  XNOR2_X1 U510 ( .A(G43GAT), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U512 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n542) );
  NAND2_X1 U514 ( .A1(n456), .A2(n542), .ZN(n458) );
  INV_X1 U515 ( .A(n571), .ZN(n464) );
  NOR2_X1 U516 ( .A1(n576), .A2(n464), .ZN(n460) );
  XNOR2_X1 U517 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(G1348GAT) );
  INV_X1 U519 ( .A(n560), .ZN(n546) );
  NOR2_X1 U520 ( .A1(n546), .A2(n464), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NOR2_X1 U524 ( .A1(n553), .A2(n464), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  NOR2_X1 U527 ( .A1(n542), .A2(n479), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT26), .B(n469), .ZN(n574) );
  AND2_X1 U529 ( .A1(n478), .A2(n574), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT95), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n542), .A2(n531), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n479), .A2(n471), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n472), .Z(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT96), .ZN(n483) );
  NAND2_X1 U537 ( .A1(n529), .A2(n478), .ZN(n538) );
  NOR2_X1 U538 ( .A1(n542), .A2(n538), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT28), .B(n479), .Z(n541) );
  INV_X1 U540 ( .A(n541), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n492), .A2(n587), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n584), .A2(n485), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n486), .Z(n528) );
  NAND2_X1 U546 ( .A1(n558), .A2(n370), .ZN(n495) );
  NOR2_X1 U547 ( .A1(n528), .A2(n495), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n511) );
  NAND2_X1 U550 ( .A1(n542), .A2(n511), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n498) );
  NAND2_X1 U552 ( .A1(n565), .A2(n553), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n491), .Z(n494) );
  NAND2_X1 U554 ( .A1(n494), .A2(n493), .ZN(n514) );
  NOR2_X1 U555 ( .A1(n495), .A2(n514), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT98), .B(n496), .ZN(n503) );
  NAND2_X1 U557 ( .A1(n529), .A2(n503), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U560 ( .A1(n503), .A2(n531), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U563 ( .A1(n503), .A2(n542), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n541), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT100), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n511), .A2(n529), .ZN(n509) );
  XOR2_X1 U569 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n507) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NAND2_X1 U573 ( .A1(n531), .A2(n511), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n513) );
  NAND2_X1 U576 ( .A1(n511), .A2(n541), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n517) );
  NAND2_X1 U579 ( .A1(n576), .A2(n560), .ZN(n527) );
  NOR2_X1 U580 ( .A1(n514), .A2(n527), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT105), .B(n515), .Z(n522) );
  NAND2_X1 U582 ( .A1(n529), .A2(n522), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n531), .A2(n522), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n519), .ZN(G1333GAT) );
  XOR2_X1 U587 ( .A(G71GAT), .B(KEYINPUT107), .Z(n521) );
  NAND2_X1 U588 ( .A1(n522), .A2(n542), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n541), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n526) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT109), .Z(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n529), .A2(n534), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n531), .A2(n534), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n542), .A2(n534), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n533), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n541), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U605 ( .A(G106GAT), .B(n537), .Z(G1339GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(n540), .Z(n556) );
  NOR2_X1 U608 ( .A1(n556), .A2(n541), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n576), .A2(n552), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1340GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n552), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  INV_X1 U616 ( .A(n552), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n549), .A2(n570), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  INV_X1 U623 ( .A(n574), .ZN(n557) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n558), .A2(n567), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XNOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n564) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT118), .Z(n562) );
  NAND2_X1 U629 ( .A1(n567), .A2(n560), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n567), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n576), .A2(n586), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n586), .A2(n370), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

