

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n551) );
  NOR2_X1 U325 ( .A1(n453), .A2(n452), .ZN(n467) );
  AND2_X1 U326 ( .A1(n558), .A2(n557), .ZN(n569) );
  XOR2_X1 U327 ( .A(n436), .B(n435), .Z(n292) );
  XOR2_X1 U328 ( .A(n404), .B(KEYINPUT21), .Z(n293) );
  XOR2_X1 U329 ( .A(n427), .B(KEYINPUT93), .Z(n294) );
  AND2_X1 U330 ( .A1(n573), .A2(n447), .ZN(n448) );
  XNOR2_X1 U331 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n403) );
  XNOR2_X1 U332 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n301) );
  XNOR2_X1 U333 ( .A(n437), .B(n292), .ZN(n438) );
  XNOR2_X1 U334 ( .A(n343), .B(n301), .ZN(n304) );
  XNOR2_X1 U335 ( .A(n439), .B(n438), .ZN(n555) );
  XNOR2_X1 U336 ( .A(n305), .B(n430), .ZN(n306) );
  XNOR2_X1 U337 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U338 ( .A1(n588), .A2(n469), .ZN(n470) );
  XNOR2_X1 U339 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U340 ( .A(n327), .B(n326), .Z(n559) );
  XOR2_X1 U341 ( .A(n425), .B(n424), .Z(n557) );
  XNOR2_X1 U342 ( .A(n472), .B(KEYINPUT38), .ZN(n481) );
  XOR2_X1 U343 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n457) );
  INV_X1 U344 ( .A(G85GAT), .ZN(n295) );
  NAND2_X1 U345 ( .A1(G92GAT), .A2(n295), .ZN(n298) );
  INV_X1 U346 ( .A(G92GAT), .ZN(n296) );
  NAND2_X1 U347 ( .A1(n296), .A2(G85GAT), .ZN(n297) );
  NAND2_X1 U348 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n343) );
  XNOR2_X1 U351 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n302) );
  XOR2_X1 U352 ( .A(G176GAT), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U353 ( .A(n302), .B(n399), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n307) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n411) );
  XOR2_X1 U356 ( .A(G57GAT), .B(KEYINPUT13), .Z(n346) );
  XNOR2_X1 U357 ( .A(n411), .B(n346), .ZN(n305) );
  XOR2_X1 U358 ( .A(G148GAT), .B(G78GAT), .Z(n430) );
  AND2_X1 U359 ( .A1(G230GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n581) );
  XOR2_X1 U361 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT74), .B(KEYINPUT76), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U364 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n313) );
  XNOR2_X1 U365 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n327) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G197GAT), .Z(n317) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(G36GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(G169GAT), .B(G8GAT), .Z(n394) );
  XOR2_X1 U372 ( .A(n318), .B(n394), .Z(n325) );
  XOR2_X1 U373 ( .A(G29GAT), .B(G43GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n335) );
  XOR2_X1 U376 ( .A(G141GAT), .B(G22GAT), .Z(n436) );
  XOR2_X1 U377 ( .A(n335), .B(n436), .Z(n322) );
  NAND2_X1 U378 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U380 ( .A(G113GAT), .B(G1GAT), .Z(n381) );
  XNOR2_X1 U381 ( .A(n323), .B(n381), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  NAND2_X1 U383 ( .A1(n581), .A2(n559), .ZN(n471) );
  XOR2_X1 U384 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n366) );
  XOR2_X1 U385 ( .A(G50GAT), .B(G162GAT), .Z(n429) );
  XOR2_X1 U386 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n329) );
  XNOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n429), .B(n330), .Z(n332) );
  NAND2_X1 U390 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n334) );
  INV_X1 U392 ( .A(KEYINPUT77), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n335), .B(KEYINPUT11), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT9), .B(KEYINPUT67), .Z(n339) );
  XNOR2_X1 U397 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U400 ( .A(G36GAT), .B(G190GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n342), .B(G218GAT), .ZN(n395) );
  XNOR2_X1 U402 ( .A(n343), .B(n395), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n546) );
  XNOR2_X1 U404 ( .A(KEYINPUT80), .B(n546), .ZN(n570) );
  INV_X1 U405 ( .A(n570), .ZN(n364) );
  XOR2_X1 U406 ( .A(n346), .B(G78GAT), .Z(n348) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G127GAT), .Z(n415) );
  XNOR2_X1 U408 ( .A(n415), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U410 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n350) );
  XNOR2_X1 U411 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U413 ( .A(n352), .B(n351), .Z(n354) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U416 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n356) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U419 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U420 ( .A(G71GAT), .B(G183GAT), .Z(n360) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G8GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n361), .B(KEYINPUT82), .ZN(n362) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n566) );
  NAND2_X1 U425 ( .A1(n364), .A2(n566), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n455) );
  XOR2_X1 U427 ( .A(KEYINPUT98), .B(KEYINPUT6), .Z(n368) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(KEYINPUT1), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U430 ( .A(G57GAT), .B(KEYINPUT5), .Z(n370) );
  XNOR2_X1 U431 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U433 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U434 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n374) );
  NAND2_X1 U435 ( .A1(G225GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U437 ( .A(KEYINPUT97), .B(n375), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U439 ( .A(G148GAT), .B(G162GAT), .Z(n379) );
  XNOR2_X1 U440 ( .A(G141GAT), .B(G127GAT), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U442 ( .A(n380), .B(G85GAT), .Z(n383) );
  XNOR2_X1 U443 ( .A(G29GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U445 ( .A(n385), .B(n384), .Z(n390) );
  XNOR2_X1 U446 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n386), .B(KEYINPUT85), .ZN(n414) );
  XOR2_X1 U448 ( .A(G155GAT), .B(KEYINPUT2), .Z(n388) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(KEYINPUT92), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n426) );
  XNOR2_X1 U451 ( .A(n414), .B(n426), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n554) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n392) );
  XNOR2_X1 U454 ( .A(KEYINPUT88), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U456 ( .A(KEYINPUT18), .B(n393), .Z(n423) );
  XOR2_X1 U457 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U460 ( .A(n398), .B(KEYINPUT99), .Z(n401) );
  XNOR2_X1 U461 ( .A(n399), .B(G92GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n423), .B(n402), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT90), .ZN(n404) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(G204GAT), .ZN(n405) );
  XOR2_X1 U466 ( .A(n293), .B(n405), .Z(n427) );
  INV_X1 U467 ( .A(n427), .ZN(n406) );
  XOR2_X2 U468 ( .A(n407), .B(n406), .Z(n550) );
  XNOR2_X1 U469 ( .A(KEYINPUT27), .B(n550), .ZN(n447) );
  NAND2_X1 U470 ( .A1(n554), .A2(n447), .ZN(n506) );
  XOR2_X1 U471 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n409) );
  XNOR2_X1 U472 ( .A(G190GAT), .B(KEYINPUT87), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U474 ( .A(n410), .B(G99GAT), .Z(n413) );
  XNOR2_X1 U475 ( .A(G43GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U477 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U478 ( .A1(G227GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U480 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U481 ( .A(G176GAT), .B(KEYINPUT89), .Z(n421) );
  XNOR2_X1 U482 ( .A(G169GAT), .B(G113GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U485 ( .A(n557), .ZN(n441) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U487 ( .A(n428), .B(n294), .ZN(n439) );
  XOR2_X1 U488 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n434) );
  XNOR2_X1 U492 ( .A(G218GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n555), .B(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n440), .B(KEYINPUT28), .ZN(n522) );
  NAND2_X1 U496 ( .A1(n441), .A2(n522), .ZN(n442) );
  NOR2_X1 U497 ( .A1(n506), .A2(n442), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n443), .B(KEYINPUT100), .ZN(n453) );
  NAND2_X1 U499 ( .A1(n557), .A2(n550), .ZN(n444) );
  NAND2_X1 U500 ( .A1(n555), .A2(n444), .ZN(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT25), .B(n445), .ZN(n450) );
  NOR2_X1 U502 ( .A1(n555), .A2(n557), .ZN(n446) );
  XNOR2_X1 U503 ( .A(KEYINPUT26), .B(n446), .ZN(n573) );
  XOR2_X1 U504 ( .A(KEYINPUT101), .B(n448), .Z(n449) );
  NOR2_X1 U505 ( .A1(n450), .A2(n449), .ZN(n451) );
  NOR2_X1 U506 ( .A1(n554), .A2(n451), .ZN(n452) );
  INV_X1 U507 ( .A(n467), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n455), .A2(n454), .ZN(n487) );
  NOR2_X1 U509 ( .A1(n471), .A2(n487), .ZN(n464) );
  NAND2_X1 U510 ( .A1(n464), .A2(n554), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U512 ( .A(G1GAT), .B(n458), .Z(G1324GAT) );
  XOR2_X1 U513 ( .A(G8GAT), .B(KEYINPUT103), .Z(n460) );
  NAND2_X1 U514 ( .A1(n464), .A2(n550), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(G1325GAT) );
  XOR2_X1 U516 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n462) );
  NAND2_X1 U517 ( .A1(n464), .A2(n557), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U519 ( .A(G15GAT), .B(n463), .ZN(G1326GAT) );
  INV_X1 U520 ( .A(n522), .ZN(n503) );
  NAND2_X1 U521 ( .A1(n503), .A2(n464), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT39), .B(KEYINPUT106), .Z(n474) );
  INV_X1 U524 ( .A(KEYINPUT36), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(n570), .ZN(n588) );
  NOR2_X1 U526 ( .A1(n467), .A2(n566), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT105), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT37), .B(n470), .ZN(n497) );
  NOR2_X1 U529 ( .A1(n471), .A2(n497), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n554), .A2(n481), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(n475), .ZN(G1328GAT) );
  NAND2_X1 U533 ( .A1(n481), .A2(n550), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U535 ( .A(G43GAT), .B(KEYINPUT107), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n478) );
  NAND2_X1 U537 ( .A1(n481), .A2(n557), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U540 ( .A(G50GAT), .B(KEYINPUT109), .Z(n483) );
  NAND2_X1 U541 ( .A1(n481), .A2(n503), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1331GAT) );
  XNOR2_X1 U543 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n489) );
  XNOR2_X1 U544 ( .A(n581), .B(KEYINPUT65), .ZN(n485) );
  INV_X1 U545 ( .A(KEYINPUT41), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n561) );
  INV_X1 U547 ( .A(n559), .ZN(n575) );
  NAND2_X1 U548 ( .A1(n561), .A2(n575), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n486), .B(KEYINPUT110), .ZN(n498) );
  NOR2_X1 U550 ( .A1(n498), .A2(n487), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n554), .A2(n493), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1332GAT) );
  NAND2_X1 U553 ( .A1(n550), .A2(n493), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U555 ( .A(G71GAT), .B(KEYINPUT111), .Z(n492) );
  NAND2_X1 U556 ( .A1(n493), .A2(n557), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n492), .B(n491), .ZN(G1334GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT43), .B(KEYINPUT112), .Z(n495) );
  NAND2_X1 U559 ( .A1(n493), .A2(n503), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G78GAT), .B(n496), .ZN(G1335GAT) );
  NOR2_X1 U562 ( .A1(n498), .A2(n497), .ZN(n502) );
  NAND2_X1 U563 ( .A1(n554), .A2(n502), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G85GAT), .B(n499), .ZN(G1336GAT) );
  NAND2_X1 U565 ( .A1(n550), .A2(n502), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U567 ( .A1(n557), .A2(n502), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U569 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT44), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G106GAT), .B(n505), .ZN(G1339GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n525) );
  INV_X1 U573 ( .A(n506), .ZN(n520) );
  AND2_X1 U574 ( .A1(n559), .A2(n561), .ZN(n508) );
  XNOR2_X1 U575 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(n510) );
  NOR2_X1 U577 ( .A1(n566), .A2(n546), .ZN(n509) );
  AND2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(KEYINPUT47), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT68), .B(KEYINPUT45), .Z(n513) );
  INV_X1 U581 ( .A(n566), .ZN(n584) );
  NOR2_X1 U582 ( .A1(n584), .A2(n588), .ZN(n512) );
  XNOR2_X1 U583 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U584 ( .A1(n559), .A2(n514), .ZN(n515) );
  NAND2_X1 U585 ( .A1(n515), .A2(n581), .ZN(n516) );
  NAND2_X1 U586 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U587 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(n549) );
  NAND2_X1 U589 ( .A1(n520), .A2(n549), .ZN(n521) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(n521), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n522), .A2(n557), .ZN(n523) );
  NOR2_X1 U592 ( .A1(n537), .A2(n523), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n534), .A2(n559), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U597 ( .A1(n534), .A2(n561), .ZN(n527) );
  XNOR2_X1 U598 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n530) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n529) );
  XNOR2_X1 U601 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(n531), .Z(n533) );
  NAND2_X1 U603 ( .A1(n534), .A2(n566), .ZN(n532) );
  XNOR2_X1 U604 ( .A(n533), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U606 ( .A1(n534), .A2(n570), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  INV_X1 U608 ( .A(n573), .ZN(n538) );
  NOR2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(KEYINPUT120), .B(n539), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n559), .A2(n547), .ZN(n540) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  NAND2_X1 U614 ( .A1(n547), .A2(n561), .ZN(n541) );
  XNOR2_X1 U615 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT121), .Z(n545) );
  NAND2_X1 U618 ( .A1(n547), .A2(n566), .ZN(n544) );
  XNOR2_X1 U619 ( .A(n545), .B(n544), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U621 ( .A(n548), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n550), .A2(n549), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n574) );
  NAND2_X1 U624 ( .A1(n555), .A2(n574), .ZN(n556) );
  XNOR2_X1 U625 ( .A(KEYINPUT55), .B(n556), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n569), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .Z(n563) );
  NAND2_X1 U629 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n569), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n575), .A2(n587), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

