//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n209), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT75), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(KEYINPUT2), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n223), .A3(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT81), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n215), .A2(new_n227), .A3(KEYINPUT2), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n215), .ZN(new_n230));
  AND2_X1   g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n233), .B2(new_n223), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n214), .B(new_n222), .C1(new_n229), .C2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n222), .B1(new_n229), .B2(new_n234), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n240));
  AND2_X1   g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n209), .B(new_n210), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT29), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n239), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n238), .A2(new_n240), .A3(new_n241), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n212), .A2(new_n236), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n214), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n243), .A2(KEYINPUT83), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n239), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(new_n238), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n203), .B(new_n245), .C1(new_n251), .C2(new_n241), .ZN(new_n252));
  INV_X1    g051(.A(new_n245), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n241), .B1(new_n250), .B2(new_n238), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n202), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G22gat), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n252), .B2(new_n255), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G64gat), .ZN(new_n263));
  INV_X1    g062(.A(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT77), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT38), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR3_X1   g073(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(KEYINPUT68), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n280), .A3(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G183gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n285), .A3(new_n273), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n288), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT28), .A3(new_n273), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT67), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n282), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n277), .B1(new_n295), .B2(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n297), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT64), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n277), .ZN(new_n303));
  NOR2_X1   g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(G190gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n313), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n302), .A4(new_n277), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n310), .A2(new_n311), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n271), .B1(new_n294), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n282), .A2(new_n289), .A3(new_n293), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n300), .A2(new_n277), .A3(new_n302), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n326), .A2(KEYINPUT64), .B1(new_n306), .B2(new_n308), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n327), .B2(new_n303), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n316), .A2(new_n313), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n307), .B(KEYINPUT65), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n320), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n325), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n271), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n236), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n270), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n213), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n310), .A2(new_n311), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n321), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n341), .B2(new_n325), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n213), .B(new_n323), .C1(new_n342), .C2(new_n271), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT37), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT87), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g144(.A(KEYINPUT76), .B(new_n270), .C1(new_n341), .C2(new_n325), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n333), .B1(new_n332), .B2(new_n271), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n213), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n343), .A2(KEYINPUT37), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n269), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n349), .A3(new_n323), .ZN(new_n355));
  XOR2_X1   g154(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n356));
  AOI21_X1  g155(.A(new_n271), .B1(new_n332), .B2(new_n236), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n324), .B2(new_n334), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n355), .B(new_n356), .C1(new_n358), .C2(new_n349), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n348), .A2(new_n213), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(KEYINPUT89), .A3(new_n355), .A4(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n270), .B1(new_n341), .B2(new_n325), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n357), .A2(new_n213), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n348), .B2(new_n213), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n265), .ZN(new_n369));
  INV_X1    g168(.A(G134gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G127gat), .ZN(new_n371));
  INV_X1    g170(.A(G127gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(KEYINPUT1), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G120gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n382), .B2(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(new_n373), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n376), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT4), .B1(new_n239), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT69), .B(G120gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n388), .B2(new_n377), .ZN(new_n389));
  INV_X1    g188(.A(new_n385), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n377), .A2(G120gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n379), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n389), .A2(new_n390), .B1(new_n392), .B2(new_n374), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n221), .A2(KEYINPUT80), .B1(new_n215), .B2(new_n218), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n233), .A2(new_n223), .B1(KEYINPUT81), .B2(new_n225), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n228), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n393), .A2(new_n396), .A3(new_n397), .A4(new_n222), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n387), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(new_n396), .A3(new_n222), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n240), .A2(new_n386), .A3(new_n235), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n239), .A2(new_n386), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n402), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n235), .A2(new_n386), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n240), .A2(new_n411), .B1(new_n387), .B2(new_n398), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G57gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G85gat), .ZN(new_n419));
  INV_X1    g218(.A(G57gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n417), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G85gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT90), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n427), .A3(new_n414), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n419), .A2(new_n423), .A3(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n405), .A2(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n428), .B(new_n429), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n436), .A3(KEYINPUT6), .A4(new_n424), .ZN(new_n437));
  AND4_X1   g236(.A1(new_n369), .A2(new_n426), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n365), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n362), .A2(new_n355), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n265), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n268), .B1(new_n364), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n261), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n369), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n358), .A2(new_n349), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT78), .B(new_n267), .C1(new_n446), .C2(new_n367), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n265), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n368), .B2(new_n266), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT85), .B1(new_n412), .B2(new_n401), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n399), .A2(new_n404), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n402), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT39), .B1(new_n408), .B2(new_n402), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n433), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT39), .B1(new_n453), .B2(new_n456), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n452), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT40), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n452), .B(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n433), .A2(new_n434), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AND4_X1   g265(.A1(new_n451), .A2(new_n462), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT82), .B1(new_n434), .B2(new_n427), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT6), .B1(new_n434), .B2(new_n427), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n415), .A2(new_n470), .A3(new_n424), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n425), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n445), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n447), .A3(new_n448), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT79), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n450), .A2(new_n447), .A3(new_n448), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g278(.A1(new_n443), .A2(new_n467), .B1(new_n261), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n393), .B1(new_n294), .B2(new_n322), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n341), .A2(new_n386), .A3(new_n325), .ZN(new_n486));
  INV_X1    g285(.A(G227gat), .ZN(new_n487));
  INV_X1    g286(.A(G233gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT32), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n490), .B2(KEYINPUT32), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT71), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n490), .B(KEYINPUT32), .C1(new_n491), .C2(new_n484), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n485), .A2(new_n486), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT72), .B1(new_n503), .B2(new_n489), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT34), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n481), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n501), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n498), .B2(new_n499), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n509), .A2(KEYINPUT74), .A3(new_n505), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n505), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT73), .B1(new_n509), .B2(new_n505), .ZN(new_n512));
  OAI22_X1  g311(.A1(new_n507), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n502), .B2(new_n506), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n505), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n509), .A2(new_n505), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(KEYINPUT36), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n480), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(new_n260), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n479), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n481), .A3(new_n506), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT74), .B1(new_n509), .B2(new_n505), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n517), .A2(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n426), .A2(new_n435), .A3(new_n437), .ZN(new_n529));
  NOR4_X1   g328(.A1(new_n260), .A2(new_n451), .A3(KEYINPUT35), .A4(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n525), .A2(KEYINPUT35), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT91), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n443), .ZN(new_n533));
  INV_X1    g332(.A(new_n467), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n479), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n260), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n526), .A2(new_n527), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT36), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n514), .B(new_n520), .C1(new_n517), .C2(new_n518), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n535), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n521), .B(new_n261), .C1(new_n511), .C2(new_n512), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT35), .B1(new_n542), .B2(new_n536), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n530), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  INV_X1    g348(.A(G1gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT16), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n549), .B2(G1gat), .ZN(new_n555));
  OAI21_X1  g354(.A(G8gat), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G15gat), .B(G22gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  INV_X1    g357(.A(G8gat), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n554), .A3(new_n559), .A4(new_n552), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G29gat), .A2(G36gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(KEYINPUT14), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n565));
  INV_X1    g364(.A(G29gat), .ZN(new_n566));
  INV_X1    g365(.A(G36gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n563), .A2(KEYINPUT14), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(G43gat), .A2(G50gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(G43gat), .A2(G50gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n572), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n570), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n568), .A2(KEYINPUT14), .A3(new_n563), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n563), .A2(KEYINPUT14), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n577), .A4(new_n562), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n562), .A4(new_n574), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n578), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n556), .A2(new_n560), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n586), .B1(new_n584), .B2(new_n578), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n548), .B(new_n585), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n548), .B(KEYINPUT13), .Z(new_n594));
  AOI21_X1  g393(.A(new_n561), .B1(new_n578), .B2(new_n584), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n585), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g396(.A(KEYINPUT96), .B(new_n561), .C1(new_n578), .C2(new_n584), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n578), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT17), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n588), .A3(new_n587), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n602), .A2(KEYINPUT18), .A3(new_n548), .A4(new_n585), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n593), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G141gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G113gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n377), .A2(G141gat), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT11), .ZN(new_n609));
  INV_X1    g408(.A(G169gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT11), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n610), .B1(new_n609), .B2(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(G197gat), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n613), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  OAI21_X1  g419(.A(G169gat), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(G197gat), .B1(new_n621), .B2(new_n614), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT92), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(G197gat), .A3(new_n614), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n623), .A2(new_n627), .A3(KEYINPUT12), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT12), .B1(new_n623), .B2(new_n627), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n604), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n632), .A2(new_n593), .A3(new_n599), .A4(new_n603), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n532), .A2(new_n547), .A3(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(G57gat), .A2(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(G57gat), .A2(G64gat), .ZN(new_n637));
  AND2_X1   g436(.A1(G71gat), .A2(G78gat), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(KEYINPUT9), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n640));
  NOR2_X1   g439(.A1(G71gat), .A2(G78gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n639), .A3(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g444(.A1(G99gat), .A2(G106gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT8), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G99gat), .B(G106gat), .ZN(new_n651));
  OAI21_X1  g450(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n652));
  AND2_X1   g451(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT7), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(new_n422), .A3(G92gat), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n650), .B(new_n651), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n422), .ZN(new_n659));
  NAND2_X1  g458(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(G92gat), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n651), .B1(new_n663), .B2(new_n650), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n643), .B(new_n645), .C1(new_n658), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n667));
  INV_X1    g466(.A(new_n651), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n644), .A2(new_n639), .A3(KEYINPUT97), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n644), .B1(new_n639), .B2(KEYINPUT97), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n669), .B(new_n657), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n665), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n665), .A2(new_n672), .A3(new_n675), .A4(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT104), .B1(new_n672), .B2(new_n666), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n658), .A2(new_n664), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n643), .A2(new_n645), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT10), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n674), .A2(new_n676), .B1(new_n678), .B2(new_n682), .ZN(new_n688));
  INV_X1    g487(.A(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT105), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n665), .A2(new_n672), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G176gat), .ZN(new_n696));
  INV_X1    g495(.A(G204gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n686), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n693), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n561), .B1(KEYINPUT21), .B2(new_n681), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n272), .ZN(new_n706));
  XNOR2_X1  g505(.A(G127gat), .B(G155gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  NAND2_X1  g507(.A1(G231gat), .A2(G233gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT98), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n708), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n706), .B(new_n711), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n681), .A2(KEYINPUT21), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n206), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n712), .B(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n600), .A2(new_n658), .A3(new_n664), .ZN(new_n718));
  NAND2_X1  g517(.A1(G232gat), .A2(G233gat), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT100), .Z(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(KEYINPUT41), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(G190gat), .B(G218gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n601), .B(new_n587), .C1(new_n658), .C2(new_n664), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n722), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n721), .A2(KEYINPUT41), .ZN(new_n728));
  XNOR2_X1  g527(.A(G134gat), .B(G162gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n726), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(new_n734), .C1(new_n726), .C2(new_n727), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n704), .A2(new_n717), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n635), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n473), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n550), .ZN(G1324gat));
  INV_X1    g540(.A(new_n739), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT16), .B(G8gat), .Z(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n451), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n451), .A4(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(new_n451), .ZN(new_n748));
  OAI21_X1  g547(.A(G8gat), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(G1325gat));
  OAI21_X1  g549(.A(new_n522), .B1(KEYINPUT36), .B2(new_n528), .ZN(new_n751));
  OAI21_X1  g550(.A(G15gat), .B1(new_n739), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n513), .A2(G15gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n739), .B2(new_n753), .ZN(G1326gat));
  NAND2_X1  g553(.A1(new_n742), .A2(new_n260), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT43), .B(G22gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1327gat));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n758));
  INV_X1    g557(.A(new_n717), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n704), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n736), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n635), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n473), .A2(G29gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n635), .A2(KEYINPUT45), .A3(new_n761), .A4(new_n763), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n736), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n532), .A2(new_n547), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n480), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n751), .A2(new_n770), .B1(new_n543), .B2(new_n544), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n771), .B2(new_n736), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n473), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n634), .A2(KEYINPUT106), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n631), .B2(new_n633), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n765), .B(new_n766), .C1(new_n780), .C2(new_n566), .ZN(G1328gat));
  NOR2_X1   g580(.A1(new_n748), .A2(G36gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT46), .B1(new_n762), .B2(new_n783), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n451), .A3(new_n772), .A4(new_n779), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G36gat), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n784), .B(new_n785), .C1(new_n789), .C2(new_n790), .ZN(G1329gat));
  INV_X1    g590(.A(new_n751), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n769), .A2(new_n792), .A3(new_n772), .A4(new_n779), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G43gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n513), .A2(G43gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n635), .A2(new_n761), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1330gat));
  NAND4_X1  g600(.A1(new_n769), .A2(new_n260), .A3(new_n772), .A4(new_n779), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G50gat), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n261), .A2(G50gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n635), .A2(new_n761), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT48), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n805), .A3(KEYINPUT48), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1331gat));
  NAND2_X1  g609(.A1(new_n541), .A2(new_n545), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n778), .A2(new_n717), .A3(new_n736), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n704), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n473), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(new_n420), .ZN(G1332gat));
  NAND2_X1  g615(.A1(new_n814), .A2(KEYINPUT108), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n818), .A3(new_n813), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n451), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT49), .B(G64gat), .Z(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(G1333gat));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n792), .A3(new_n819), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G71gat), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n814), .A2(G71gat), .A3(new_n513), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(KEYINPUT50), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1334gat));
  NAND2_X1  g631(.A1(new_n820), .A2(new_n260), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT109), .B(G78gat), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(G1335gat));
  NOR2_X1   g634(.A1(new_n775), .A2(new_n777), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n717), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n704), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n773), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G85gat), .B1(new_n840), .B2(new_n473), .ZN(new_n841));
  INV_X1    g640(.A(new_n736), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n842), .A3(new_n837), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(new_n422), .A3(new_n774), .A4(new_n703), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(G1336gat));
  NAND4_X1  g646(.A1(new_n769), .A2(new_n451), .A3(new_n772), .A4(new_n839), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G92gat), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n703), .A2(new_n264), .A3(new_n451), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT110), .Z(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n849), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n849), .B(new_n858), .C1(new_n852), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1337gat));
  OAI21_X1  g659(.A(G99gat), .B1(new_n840), .B2(new_n751), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n513), .A2(G99gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n703), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1338gat));
  NOR3_X1   g663(.A1(new_n704), .A2(new_n261), .A3(G106gat), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT111), .Z(new_n866));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n845), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n769), .A2(new_n260), .A3(new_n772), .A4(new_n839), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G106gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n868), .A2(new_n869), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n866), .B1(new_n850), .B2(new_n851), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(G106gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n877), .ZN(G1339gat));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n687), .A2(new_n690), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n688), .A2(new_n689), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n701), .A2(KEYINPUT54), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT55), .A4(new_n699), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n684), .B2(new_n686), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n881), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(KEYINPUT114), .A3(new_n699), .A4(new_n880), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n702), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n880), .A2(new_n699), .A3(new_n882), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n836), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n597), .A2(new_n598), .A3(new_n594), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n548), .B1(new_n602), .B2(new_n585), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n896), .A2(new_n897), .B1(new_n618), .B2(new_n622), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n633), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n700), .B2(new_n702), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n894), .B2(new_n901), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n842), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n736), .A2(new_n899), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n906), .A3(new_n893), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n759), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n812), .A2(new_n703), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n260), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n520), .B1(new_n517), .B2(new_n518), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n451), .A2(new_n473), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G113gat), .B1(new_n917), .B2(new_n836), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n513), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n377), .B1(new_n631), .B2(new_n633), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(G1340gat));
  OAI21_X1  g723(.A(G120gat), .B1(new_n921), .B2(new_n704), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n703), .A2(new_n382), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n916), .B2(new_n926), .ZN(G1341gat));
  OAI21_X1  g726(.A(G127gat), .B1(new_n921), .B2(new_n759), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n717), .A2(new_n372), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n916), .B2(new_n929), .ZN(G1342gat));
  NAND2_X1  g729(.A1(new_n842), .A2(new_n370), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n916), .A2(KEYINPUT56), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G134gat), .B1(new_n921), .B2(new_n736), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT56), .B1(new_n916), .B2(new_n931), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G1343gat));
  NOR2_X1   g734(.A1(new_n792), .A2(new_n919), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n894), .A2(new_n901), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n842), .B1(new_n937), .B2(KEYINPUT115), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n908), .B1(new_n938), .B2(new_n902), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n912), .B1(new_n939), .B2(new_n717), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n940), .B2(new_n260), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n261), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n634), .A2(new_n702), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n892), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n900), .B1(new_n947), .B2(new_n890), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n907), .B1(new_n948), .B2(new_n842), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n759), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n944), .B1(new_n912), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n634), .B(new_n936), .C1(new_n941), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G141gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n940), .A2(new_n260), .ZN(new_n954));
  INV_X1    g753(.A(new_n936), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n634), .A2(new_n605), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(KEYINPUT58), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT58), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n836), .B(new_n936), .C1(new_n941), .C2(new_n951), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(G141gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(G1344gat));
  AOI21_X1  g762(.A(new_n261), .B1(new_n909), .B2(new_n912), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n936), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n704), .A2(G148gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(KEYINPUT117), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT117), .ZN(new_n969));
  INV_X1    g768(.A(new_n967), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT59), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G148gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n942), .ZN(new_n975));
  INV_X1    g774(.A(new_n951), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n955), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n977), .B2(new_n703), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n737), .A2(new_n634), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n979), .B1(new_n949), .B2(new_n759), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n942), .B1(new_n980), .B2(new_n261), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT118), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(KEYINPUT118), .B(new_n942), .C1(new_n980), .C2(new_n261), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n944), .B1(new_n909), .B2(new_n912), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n703), .B(new_n936), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n973), .B1(new_n987), .B2(G148gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n972), .B1(new_n978), .B2(new_n988), .ZN(G1345gat));
  NAND4_X1  g788(.A1(new_n940), .A2(new_n260), .A3(new_n717), .A4(new_n936), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n216), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n936), .B1(new_n941), .B2(new_n951), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n717), .A2(G155gat), .ZN(new_n993));
  XOR2_X1   g792(.A(new_n993), .B(KEYINPUT119), .Z(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT120), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g796(.A(KEYINPUT120), .B(new_n991), .C1(new_n992), .C2(new_n994), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(G1346gat));
  OAI21_X1  g798(.A(G162gat), .B1(new_n992), .B2(new_n736), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n966), .A2(new_n217), .A3(new_n842), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1347gat));
  NAND2_X1  g801(.A1(new_n451), .A2(new_n473), .ZN(new_n1003));
  INV_X1    g802(.A(new_n1003), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n913), .A2(new_n914), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(G169gat), .B1(new_n1005), .B2(new_n836), .ZN(new_n1006));
  XOR2_X1   g805(.A(new_n1003), .B(KEYINPUT121), .Z(new_n1007));
  NOR2_X1   g806(.A1(new_n1007), .A2(new_n513), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n913), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n610), .B1(new_n631), .B2(new_n633), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(G1348gat));
  INV_X1    g811(.A(G176gat), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1005), .A2(new_n1013), .A3(new_n703), .ZN(new_n1014));
  OAI21_X1  g813(.A(G176gat), .B1(new_n1009), .B2(new_n704), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(G1349gat));
  NAND4_X1  g815(.A1(new_n940), .A2(new_n261), .A3(new_n717), .A4(new_n1008), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT123), .ZN(new_n1018));
  AOI22_X1  g817(.A1(new_n1017), .A2(G183gat), .B1(new_n1018), .B2(KEYINPUT60), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n717), .A2(new_n291), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n913), .A2(new_n914), .A3(new_n1004), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT122), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1018), .B1(new_n1022), .B2(KEYINPUT60), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT124), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1024), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1026));
  NOR2_X1   g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1350gat));
  NAND4_X1  g826(.A1(new_n940), .A2(new_n261), .A3(new_n842), .A4(new_n1008), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1028), .A2(G190gat), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1029), .A2(KEYINPUT125), .ZN(new_n1030));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1028), .A2(new_n1031), .A3(G190gat), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1005), .A2(new_n273), .A3(new_n842), .ZN(new_n1034));
  OAI211_X1 g833(.A(new_n1033), .B(new_n1034), .C1(KEYINPUT61), .C2(new_n1030), .ZN(G1351gat));
  NOR2_X1   g834(.A1(new_n261), .A2(new_n748), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n751), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n751), .A2(KEYINPUT126), .A3(new_n1036), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n774), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AND2_X1   g840(.A1(new_n1041), .A2(new_n940), .ZN(new_n1042));
  AOI21_X1  g841(.A(G197gat), .B1(new_n1042), .B2(new_n836), .ZN(new_n1043));
  NOR2_X1   g842(.A1(new_n985), .A2(new_n986), .ZN(new_n1044));
  NOR3_X1   g843(.A1(new_n1044), .A2(new_n792), .A3(new_n1007), .ZN(new_n1045));
  AOI21_X1  g844(.A(new_n617), .B1(new_n631), .B2(new_n633), .ZN(new_n1046));
  AOI21_X1  g845(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G1352gat));
  NOR2_X1   g846(.A1(new_n792), .A2(new_n1007), .ZN(new_n1048));
  OAI211_X1 g847(.A(new_n703), .B(new_n1048), .C1(new_n985), .C2(new_n986), .ZN(new_n1049));
  NAND2_X1  g848(.A1(new_n1049), .A2(G204gat), .ZN(new_n1050));
  NAND4_X1  g849(.A1(new_n1041), .A2(new_n697), .A3(new_n703), .A4(new_n940), .ZN(new_n1051));
  NAND2_X1  g850(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1052));
  OR2_X1    g851(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1053));
  NAND3_X1  g852(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(G1353gat));
  NAND3_X1  g853(.A1(new_n1042), .A2(new_n206), .A3(new_n717), .ZN(new_n1055));
  OAI211_X1 g854(.A(new_n717), .B(new_n1048), .C1(new_n985), .C2(new_n986), .ZN(new_n1056));
  AND3_X1   g855(.A1(new_n1056), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1057));
  AOI21_X1  g856(.A(KEYINPUT63), .B1(new_n1056), .B2(G211gat), .ZN(new_n1058));
  OAI21_X1  g857(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(G1354gat));
  AOI21_X1  g858(.A(G218gat), .B1(new_n1042), .B2(new_n842), .ZN(new_n1060));
  NOR2_X1   g859(.A1(new_n736), .A2(new_n207), .ZN(new_n1061));
  AOI21_X1  g860(.A(new_n1060), .B1(new_n1045), .B2(new_n1061), .ZN(G1355gat));
endmodule


