

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580;

  XOR2_X1 U318 ( .A(G99GAT), .B(KEYINPUT69), .Z(n286) );
  XNOR2_X1 U319 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n368) );
  XNOR2_X1 U320 ( .A(n369), .B(n368), .ZN(n370) );
  AND2_X1 U321 ( .A1(n505), .A2(n405), .ZN(n562) );
  XNOR2_X1 U322 ( .A(n377), .B(n376), .ZN(n569) );
  XNOR2_X1 U323 ( .A(n443), .B(G183GAT), .ZN(n444) );
  XNOR2_X1 U324 ( .A(n445), .B(n444), .ZN(G1350GAT) );
  XOR2_X1 U325 ( .A(G22GAT), .B(G78GAT), .Z(n288) );
  XOR2_X1 U326 ( .A(G57GAT), .B(KEYINPUT13), .Z(n373) );
  XOR2_X1 U327 ( .A(G183GAT), .B(G8GAT), .Z(n400) );
  XNOR2_X1 U328 ( .A(n373), .B(n400), .ZN(n287) );
  XNOR2_X1 U329 ( .A(n288), .B(n287), .ZN(n289) );
  XOR2_X1 U330 ( .A(n289), .B(G71GAT), .Z(n295) );
  XNOR2_X1 U331 ( .A(G1GAT), .B(G15GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n290), .B(KEYINPUT67), .ZN(n349) );
  XOR2_X1 U333 ( .A(n349), .B(KEYINPUT76), .Z(n292) );
  NAND2_X1 U334 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n293) );
  XNOR2_X1 U336 ( .A(G127GAT), .B(n293), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n303) );
  XOR2_X1 U338 ( .A(KEYINPUT15), .B(G64GAT), .Z(n297) );
  XNOR2_X1 U339 ( .A(G155GAT), .B(G211GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U341 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n299) );
  XNOR2_X1 U342 ( .A(KEYINPUT12), .B(KEYINPUT77), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U344 ( .A(n301), .B(n300), .Z(n302) );
  XNOR2_X1 U345 ( .A(n303), .B(n302), .ZN(n573) );
  INV_X1 U346 ( .A(n573), .ZN(n545) );
  XNOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n304), .B(KEYINPUT2), .ZN(n415) );
  XOR2_X1 U349 ( .A(G85GAT), .B(n415), .Z(n306) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(G120GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U352 ( .A(G162GAT), .B(n307), .ZN(n328) );
  XOR2_X1 U353 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n309) );
  XNOR2_X1 U354 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT4), .B(n310), .Z(n312) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(n313), .B(KEYINPUT91), .Z(n318) );
  XOR2_X1 U360 ( .A(KEYINPUT78), .B(G134GAT), .Z(n315) );
  XNOR2_X1 U361 ( .A(G127GAT), .B(G113GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U363 ( .A(KEYINPUT0), .B(n316), .ZN(n440) );
  XOR2_X1 U364 ( .A(n440), .B(KEYINPUT1), .Z(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n326) );
  XOR2_X1 U366 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n320) );
  XNOR2_X1 U367 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U369 ( .A(G1GAT), .B(G57GAT), .Z(n322) );
  XNOR2_X1 U370 ( .A(G148GAT), .B(G141GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n479) );
  INV_X1 U375 ( .A(n479), .ZN(n505) );
  XOR2_X1 U376 ( .A(KEYINPUT11), .B(G92GAT), .Z(n330) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(G106GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n332) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(KEYINPUT73), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U382 ( .A(n334), .B(n333), .Z(n343) );
  XOR2_X1 U383 ( .A(KEYINPUT66), .B(KEYINPUT7), .Z(n336) );
  XNOR2_X1 U384 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(n337), .ZN(n361) );
  XOR2_X1 U387 ( .A(G190GAT), .B(G36GAT), .Z(n390) );
  XNOR2_X1 U388 ( .A(G162GAT), .B(G50GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n338), .B(KEYINPUT72), .ZN(n407) );
  XNOR2_X1 U390 ( .A(n390), .B(n407), .ZN(n340) );
  AND2_X1 U391 ( .A1(G232GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U393 ( .A(n361), .B(n341), .Z(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n345) );
  INV_X1 U395 ( .A(KEYINPUT74), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n348) );
  XNOR2_X1 U397 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n286), .B(n346), .ZN(n369) );
  XNOR2_X1 U399 ( .A(G134GAT), .B(n369), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n556) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .Z(n414) );
  XOR2_X1 U402 ( .A(n414), .B(n349), .Z(n351) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n353) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U408 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U409 ( .A(G197GAT), .B(G169GAT), .Z(n357) );
  XNOR2_X1 U410 ( .A(G113GAT), .B(G8GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n358), .B(KEYINPUT29), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n563) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  XOR2_X1 U416 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U417 ( .A(n363), .B(n431), .ZN(n377) );
  XOR2_X1 U418 ( .A(G204GAT), .B(G176GAT), .Z(n365) );
  XNOR2_X1 U419 ( .A(G92GAT), .B(G64GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n391) );
  XOR2_X1 U421 ( .A(KEYINPUT68), .B(G78GAT), .Z(n367) );
  XNOR2_X1 U422 ( .A(G148GAT), .B(G106GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n406) );
  XNOR2_X1 U424 ( .A(n391), .B(n406), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U426 ( .A(n372), .B(KEYINPUT31), .Z(n375) );
  XNOR2_X1 U427 ( .A(n373), .B(KEYINPUT33), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U429 ( .A(KEYINPUT41), .B(n569), .ZN(n553) );
  NOR2_X1 U430 ( .A1(n563), .A2(n553), .ZN(n378) );
  XOR2_X1 U431 ( .A(n378), .B(KEYINPUT46), .Z(n379) );
  NAND2_X1 U432 ( .A1(n556), .A2(n379), .ZN(n380) );
  NOR2_X1 U433 ( .A1(n573), .A2(n380), .ZN(n381) );
  XOR2_X1 U434 ( .A(n381), .B(KEYINPUT47), .Z(n388) );
  INV_X1 U435 ( .A(KEYINPUT45), .ZN(n383) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(n556), .Z(n576) );
  NAND2_X1 U437 ( .A1(n576), .A2(n573), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n563), .A2(n384), .ZN(n385) );
  NOR2_X1 U440 ( .A1(n569), .A2(n385), .ZN(n386) );
  XNOR2_X1 U441 ( .A(KEYINPUT112), .B(n386), .ZN(n387) );
  NOR2_X1 U442 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U443 ( .A(KEYINPUT48), .B(n389), .ZN(n517) );
  XOR2_X1 U444 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U447 ( .A(KEYINPUT84), .B(G197GAT), .Z(n395) );
  XNOR2_X1 U448 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U450 ( .A(G211GAT), .B(n396), .Z(n424) );
  XOR2_X1 U451 ( .A(n397), .B(n424), .Z(n402) );
  XOR2_X1 U452 ( .A(G169GAT), .B(KEYINPUT19), .Z(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n435) );
  XNOR2_X1 U455 ( .A(n400), .B(n435), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n482) );
  XNOR2_X1 U457 ( .A(KEYINPUT119), .B(n482), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n517), .A2(n403), .ZN(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT54), .B(n404), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n422) );
  XOR2_X1 U461 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n409) );
  XNOR2_X1 U462 ( .A(KEYINPUT82), .B(KEYINPUT86), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U464 ( .A(KEYINPUT85), .B(n410), .Z(n412) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U467 ( .A(n413), .B(KEYINPUT24), .Z(n420) );
  XOR2_X1 U468 ( .A(KEYINPUT83), .B(n414), .Z(n417) );
  XNOR2_X1 U469 ( .A(n415), .B(G204GAT), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n418), .B(KEYINPUT87), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(n423), .ZN(n458) );
  NAND2_X1 U475 ( .A1(n562), .A2(n458), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n425), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U477 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n427) );
  XNOR2_X1 U478 ( .A(G15GAT), .B(G176GAT), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n439) );
  XOR2_X1 U480 ( .A(G183GAT), .B(G190GAT), .Z(n429) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G99GAT), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U483 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U486 ( .A(n434), .B(KEYINPUT81), .Z(n437) );
  XNOR2_X1 U487 ( .A(n435), .B(KEYINPUT80), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U490 ( .A(n441), .B(n440), .ZN(n485) );
  NAND2_X1 U491 ( .A1(n442), .A2(n485), .ZN(n557) );
  NOR2_X1 U492 ( .A1(n545), .A2(n557), .ZN(n445) );
  XNOR2_X1 U493 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n447) );
  XNOR2_X1 U495 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n466) );
  NOR2_X1 U497 ( .A1(n563), .A2(n569), .ZN(n476) );
  NAND2_X1 U498 ( .A1(n482), .A2(n485), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n448), .B(KEYINPUT96), .ZN(n449) );
  NAND2_X1 U500 ( .A1(n449), .A2(n458), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n450), .B(KEYINPUT25), .ZN(n454) );
  XOR2_X1 U502 ( .A(n482), .B(KEYINPUT27), .Z(n459) );
  XOR2_X1 U503 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n452) );
  OR2_X1 U504 ( .A1(n458), .A2(n485), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n537) );
  NOR2_X1 U506 ( .A1(n459), .A2(n537), .ZN(n453) );
  NOR2_X1 U507 ( .A1(n454), .A2(n453), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT97), .B(n455), .Z(n456) );
  NOR2_X1 U509 ( .A1(n479), .A2(n456), .ZN(n457) );
  XNOR2_X1 U510 ( .A(KEYINPUT98), .B(n457), .ZN(n462) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT28), .ZN(n521) );
  INV_X1 U512 ( .A(n521), .ZN(n489) );
  NOR2_X1 U513 ( .A1(n505), .A2(n459), .ZN(n519) );
  INV_X1 U514 ( .A(n485), .ZN(n523) );
  NAND2_X1 U515 ( .A1(n519), .A2(n523), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n489), .A2(n460), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n473) );
  NAND2_X1 U518 ( .A1(n556), .A2(n573), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT16), .B(n463), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n473), .A2(n464), .ZN(n492) );
  NAND2_X1 U521 ( .A1(n476), .A2(n492), .ZN(n470) );
  NOR2_X1 U522 ( .A1(n505), .A2(n470), .ZN(n465) );
  XOR2_X1 U523 ( .A(n466), .B(n465), .Z(G1324GAT) );
  INV_X1 U524 ( .A(n482), .ZN(n507) );
  NOR2_X1 U525 ( .A1(n507), .A2(n470), .ZN(n467) );
  XOR2_X1 U526 ( .A(G8GAT), .B(n467), .Z(G1325GAT) );
  NOR2_X1 U527 ( .A1(n523), .A2(n470), .ZN(n469) );
  XNOR2_X1 U528 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(G1326GAT) );
  NOR2_X1 U530 ( .A1(n521), .A2(n470), .ZN(n472) );
  XNOR2_X1 U531 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(G1327GAT) );
  XOR2_X1 U533 ( .A(G29GAT), .B(KEYINPUT39), .Z(n481) );
  XOR2_X1 U534 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n478) );
  NOR2_X1 U535 ( .A1(n573), .A2(n473), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n576), .A2(n474), .ZN(n475) );
  XNOR2_X1 U537 ( .A(KEYINPUT37), .B(n475), .ZN(n504) );
  NAND2_X1 U538 ( .A1(n476), .A2(n504), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n488), .A2(n479), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(G1328GAT) );
  XOR2_X1 U542 ( .A(G36GAT), .B(KEYINPUT103), .Z(n484) );
  NAND2_X1 U543 ( .A1(n488), .A2(n482), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1329GAT) );
  NAND2_X1 U545 ( .A1(n485), .A2(n488), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT40), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G43GAT), .B(n487), .ZN(G1330GAT) );
  NAND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U550 ( .A(n563), .ZN(n524) );
  NOR2_X1 U551 ( .A1(n553), .A2(n524), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(n491), .Z(n503) );
  NAND2_X1 U553 ( .A1(n503), .A2(n492), .ZN(n500) );
  NOR2_X1 U554 ( .A1(n505), .A2(n500), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U557 ( .A(G57GAT), .B(n495), .Z(G1332GAT) );
  NOR2_X1 U558 ( .A1(n507), .A2(n500), .ZN(n496) );
  XOR2_X1 U559 ( .A(KEYINPUT106), .B(n496), .Z(n497) );
  XNOR2_X1 U560 ( .A(G64GAT), .B(n497), .ZN(G1333GAT) );
  NOR2_X1 U561 ( .A1(n523), .A2(n500), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1334GAT) );
  NOR2_X1 U564 ( .A1(n521), .A2(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  NAND2_X1 U567 ( .A1(n504), .A2(n503), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n505), .A2(n513), .ZN(n506) );
  XOR2_X1 U569 ( .A(G85GAT), .B(n506), .Z(G1336GAT) );
  NOR2_X1 U570 ( .A1(n507), .A2(n513), .ZN(n509) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G92GAT), .B(n510), .ZN(G1337GAT) );
  NOR2_X1 U574 ( .A1(n523), .A2(n513), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT110), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(G99GAT), .B(n512), .ZN(G1338GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  INV_X1 U581 ( .A(n517), .ZN(n518) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(KEYINPUT113), .B(n520), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n521), .A2(n538), .ZN(n522) );
  NOR2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n533), .A2(n524), .ZN(n525) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  INV_X1 U589 ( .A(n553), .ZN(n526) );
  NAND2_X1 U590 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  NAND2_X1 U592 ( .A1(n573), .A2(n533), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n532) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n536) );
  INV_X1 U598 ( .A(n556), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U600 ( .A(n536), .B(n535), .Z(G1343GAT) );
  INV_X1 U601 ( .A(n537), .ZN(n561) );
  NAND2_X1 U602 ( .A1(n538), .A2(n561), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n563), .A2(n547), .ZN(n539) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n539), .Z(n540) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(n540), .ZN(G1344GAT) );
  NOR2_X1 U606 ( .A1(n547), .A2(n553), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n542) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n547), .ZN(n546) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  NOR2_X1 U613 ( .A1(n556), .A2(n547), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(n548), .Z(n549) );
  XNOR2_X1 U615 ( .A(G162GAT), .B(n549), .ZN(G1347GAT) );
  NOR2_X1 U616 ( .A1(n563), .A2(n557), .ZN(n550) );
  XOR2_X1 U617 ( .A(G169GAT), .B(n550), .Z(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n552) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n557), .A2(n553), .ZN(n554) );
  XOR2_X1 U622 ( .A(n555), .B(n554), .Z(G1349GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n568) );
  NOR2_X1 U628 ( .A1(n563), .A2(n568), .ZN(n567) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT124), .B(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U634 ( .A(n568), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n577), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

