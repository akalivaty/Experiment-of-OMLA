

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  XOR2_X1 U324 ( .A(n464), .B(n425), .Z(n531) );
  XNOR2_X1 U325 ( .A(n502), .B(KEYINPUT37), .ZN(n526) );
  INV_X1 U326 ( .A(n526), .ZN(n527) );
  XOR2_X1 U327 ( .A(KEYINPUT28), .B(n476), .Z(n543) );
  XOR2_X1 U328 ( .A(KEYINPUT98), .B(n475), .Z(n292) );
  XOR2_X1 U329 ( .A(KEYINPUT92), .B(n414), .Z(n293) );
  XOR2_X1 U330 ( .A(n452), .B(n414), .Z(n294) );
  XNOR2_X1 U331 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n354) );
  XNOR2_X1 U332 ( .A(n355), .B(n354), .ZN(n370) );
  XNOR2_X1 U333 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U334 ( .A(n407), .B(n406), .ZN(n539) );
  XNOR2_X1 U335 ( .A(n294), .B(n367), .ZN(n335) );
  NOR2_X1 U336 ( .A1(n529), .A2(n429), .ZN(n584) );
  XNOR2_X1 U337 ( .A(n336), .B(n335), .ZN(n566) );
  XNOR2_X1 U338 ( .A(KEYINPUT38), .B(n505), .ZN(n513) );
  XNOR2_X1 U339 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U340 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G120GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(G29GAT), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(G57GAT), .B(G155GAT), .Z(n298) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(G148GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n302) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U351 ( .A(KEYINPUT4), .B(n303), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n314) );
  XOR2_X1 U353 ( .A(KEYINPUT89), .B(KEYINPUT91), .Z(n307) );
  XNOR2_X1 U354 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n312) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n308), .B(KEYINPUT2), .ZN(n441) );
  XOR2_X1 U358 ( .A(n441), .B(G162GAT), .Z(n310) );
  XOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .Z(n458) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(n458), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U362 ( .A(n312), .B(n311), .Z(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n529) );
  INV_X1 U364 ( .A(KEYINPUT54), .ZN(n428) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n315), .B(KEYINPUT7), .ZN(n389) );
  INV_X1 U367 ( .A(n389), .ZN(n316) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  NAND2_X1 U369 ( .A1(n316), .A2(n440), .ZN(n319) );
  INV_X1 U370 ( .A(n440), .ZN(n317) );
  NAND2_X1 U371 ( .A1(n317), .A2(n389), .ZN(n318) );
  NAND2_X1 U372 ( .A1(n319), .A2(n318), .ZN(n321) );
  NAND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n327) );
  INV_X1 U375 ( .A(n327), .ZN(n325) );
  XOR2_X1 U376 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n323) );
  XNOR2_X1 U377 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n326) );
  INV_X1 U379 ( .A(n326), .ZN(n324) );
  NAND2_X1 U380 ( .A1(n325), .A2(n324), .ZN(n329) );
  NAND2_X1 U381 ( .A1(n327), .A2(n326), .ZN(n328) );
  NAND2_X1 U382 ( .A1(n329), .A2(n328), .ZN(n336) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n330), .B(G134GAT), .ZN(n452) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G218GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n331), .B(KEYINPUT75), .ZN(n414) );
  XOR2_X1 U387 ( .A(KEYINPUT72), .B(G92GAT), .Z(n333) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(n334), .ZN(n367) );
  XOR2_X1 U391 ( .A(n566), .B(KEYINPUT76), .Z(n552) );
  XNOR2_X1 U392 ( .A(KEYINPUT36), .B(n552), .ZN(n499) );
  XOR2_X1 U393 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n338) );
  XNOR2_X1 U394 ( .A(KEYINPUT13), .B(G64GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(G57GAT), .B(n339), .Z(n366) );
  XOR2_X1 U397 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n341) );
  XNOR2_X1 U398 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n366), .B(n342), .ZN(n353) );
  XOR2_X1 U401 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n344) );
  XNOR2_X1 U402 ( .A(G71GAT), .B(G78GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(G8GAT), .B(G211GAT), .Z(n419) );
  XOR2_X1 U405 ( .A(n345), .B(n419), .Z(n351) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(G1GAT), .Z(n385) );
  XOR2_X1 U407 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XNOR2_X1 U408 ( .A(G15GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n346), .B(G127GAT), .ZN(n457) );
  XOR2_X1 U410 ( .A(n439), .B(n457), .Z(n348) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n385), .B(n349), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(n353), .B(n352), .Z(n486) );
  INV_X1 U416 ( .A(n486), .ZN(n594) );
  NAND2_X1 U417 ( .A1(n499), .A2(n594), .ZN(n355) );
  XOR2_X1 U418 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U419 ( .A(KEYINPUT70), .B(KEYINPUT33), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U421 ( .A(n358), .B(G204GAT), .Z(n360) );
  XOR2_X1 U422 ( .A(G120GAT), .B(G71GAT), .Z(n459) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(n459), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U425 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n361), .B(G148GAT), .ZN(n436) );
  XOR2_X1 U427 ( .A(n436), .B(KEYINPUT73), .Z(n363) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n395) );
  NOR2_X1 U433 ( .A1(n370), .A2(n395), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n371), .B(KEYINPUT113), .ZN(n394) );
  XOR2_X1 U435 ( .A(G141GAT), .B(G22GAT), .Z(n373) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G15GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U438 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n375) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(G8GAT), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n393) );
  INV_X1 U442 ( .A(G36GAT), .ZN(n378) );
  NAND2_X1 U443 ( .A1(G113GAT), .A2(n378), .ZN(n381) );
  INV_X1 U444 ( .A(G113GAT), .ZN(n379) );
  NAND2_X1 U445 ( .A1(n379), .A2(G36GAT), .ZN(n380) );
  NAND2_X1 U446 ( .A1(n381), .A2(n380), .ZN(n383) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(G43GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U449 ( .A(n385), .B(n384), .Z(n387) );
  NAND2_X1 U450 ( .A1(G229GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U452 ( .A(n388), .B(KEYINPUT29), .Z(n391) );
  XNOR2_X1 U453 ( .A(n389), .B(KEYINPUT66), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n585) );
  INV_X1 U456 ( .A(n585), .ZN(n558) );
  NOR2_X1 U457 ( .A1(n394), .A2(n558), .ZN(n403) );
  XOR2_X1 U458 ( .A(KEYINPUT109), .B(n594), .Z(n579) );
  XOR2_X1 U459 ( .A(KEYINPUT41), .B(n395), .Z(n560) );
  INV_X1 U460 ( .A(n560), .ZN(n576) );
  NOR2_X1 U461 ( .A1(n585), .A2(n576), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT46), .ZN(n397) );
  NOR2_X1 U463 ( .A1(n579), .A2(n397), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n398), .B(KEYINPUT110), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n399), .A2(n566), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT47), .ZN(n401) );
  XOR2_X1 U467 ( .A(n401), .B(KEYINPUT111), .Z(n402) );
  NOR2_X1 U468 ( .A1(n403), .A2(n402), .ZN(n407) );
  INV_X1 U469 ( .A(KEYINPUT48), .ZN(n405) );
  INV_X1 U470 ( .A(KEYINPUT64), .ZN(n404) );
  XOR2_X1 U471 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT17), .B(G176GAT), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U474 ( .A(G169GAT), .B(n410), .Z(n464) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n412) );
  XNOR2_X1 U476 ( .A(KEYINPUT86), .B(G204GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U478 ( .A(G197GAT), .B(n413), .Z(n448) );
  NAND2_X1 U479 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n293), .B(n415), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n448), .B(n416), .ZN(n424) );
  XOR2_X1 U482 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n418) );
  XNOR2_X1 U483 ( .A(G183GAT), .B(G64GAT), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U485 ( .A(n420), .B(n419), .Z(n422) );
  XNOR2_X1 U486 ( .A(G190GAT), .B(G92GAT), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U489 ( .A(n531), .ZN(n426) );
  NOR2_X1 U490 ( .A1(n539), .A2(n426), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n431) );
  XNOR2_X1 U493 ( .A(G218GAT), .B(G106GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n433) );
  XNOR2_X1 U496 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n446) );
  XOR2_X1 U499 ( .A(n436), .B(G211GAT), .Z(n438) );
  NAND2_X1 U500 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n476) );
  NAND2_X1 U507 ( .A1(n584), .A2(n476), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n449), .B(KEYINPUT55), .ZN(n465) );
  XOR2_X1 U509 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n451) );
  XNOR2_X1 U510 ( .A(G99GAT), .B(KEYINPUT82), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(n456) );
  XOR2_X1 U512 ( .A(n452), .B(KEYINPUT20), .Z(n454) );
  NAND2_X1 U513 ( .A1(G227GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n540) );
  NAND2_X1 U520 ( .A1(n465), .A2(n540), .ZN(n575) );
  INV_X1 U521 ( .A(n575), .ZN(n580) );
  NAND2_X1 U522 ( .A1(n580), .A2(n552), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n467) );
  INV_X1 U524 ( .A(G190GAT), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n490) );
  NOR2_X1 U526 ( .A1(n585), .A2(n395), .ZN(n503) );
  XNOR2_X1 U527 ( .A(KEYINPUT83), .B(n540), .ZN(n471) );
  XNOR2_X1 U528 ( .A(KEYINPUT27), .B(n531), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n529), .A2(n480), .ZN(n538) );
  NOR2_X1 U530 ( .A1(n543), .A2(n538), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT95), .ZN(n485) );
  NAND2_X1 U533 ( .A1(n540), .A2(n531), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n473), .A2(n476), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT25), .ZN(n475) );
  NOR2_X1 U536 ( .A1(n540), .A2(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT96), .B(n479), .Z(n583) );
  NAND2_X1 U540 ( .A1(n583), .A2(n480), .ZN(n481) );
  NAND2_X1 U541 ( .A1(n292), .A2(n481), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT99), .B(n482), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n529), .A2(n483), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n500) );
  NOR2_X1 U545 ( .A1(n486), .A2(n552), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U547 ( .A1(n500), .A2(n488), .ZN(n516) );
  AND2_X1 U548 ( .A1(n503), .A2(n516), .ZN(n497) );
  NAND2_X1 U549 ( .A1(n497), .A2(n529), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n491), .Z(G1324GAT) );
  XOR2_X1 U552 ( .A(G8GAT), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U553 ( .A1(n497), .A2(n531), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n495) );
  NAND2_X1 U556 ( .A1(n497), .A2(n540), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  NAND2_X1 U559 ( .A1(n543), .A2(n497), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n507) );
  NOR2_X1 U562 ( .A1(n594), .A2(n500), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n499), .A2(n501), .ZN(n502) );
  NAND2_X1 U564 ( .A1(n526), .A2(n503), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(KEYINPUT103), .ZN(n505) );
  NAND2_X1 U566 ( .A1(n513), .A2(n529), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n508), .ZN(G1328GAT) );
  XOR2_X1 U569 ( .A(G36GAT), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U570 ( .A1(n531), .A2(n513), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n540), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n543), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U578 ( .A1(n560), .A2(n585), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(KEYINPUT106), .ZN(n528) );
  INV_X1 U580 ( .A(n516), .ZN(n517) );
  NOR2_X1 U581 ( .A1(n528), .A2(n517), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n529), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n531), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n540), .A2(n523), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n543), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n529), .A2(n535), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n535), .A2(n531), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n540), .A2(n535), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT108), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(n534), .ZN(G1338GAT) );
  NAND2_X1 U600 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT115), .Z(n545) );
  NOR2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n556) );
  NAND2_X1 U605 ( .A1(n556), .A2(n540), .ZN(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT114), .B(n541), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n553), .A2(n558), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U611 ( .A1(n553), .A2(n560), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n550) );
  NAND2_X1 U615 ( .A1(n553), .A2(n579), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n583), .A2(n556), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(n557), .Z(n568) );
  NAND2_X1 U623 ( .A1(n558), .A2(n568), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n568), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT52), .Z(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n568), .A2(n594), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U632 ( .A(n566), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT120), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n570), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n585), .A2(n575), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n574) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(n578), .B(n577), .Z(G1349GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT123), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1350GAT) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n591) );
  NOR2_X1 U648 ( .A1(n585), .A2(n591), .ZN(n590) );
  XOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n587) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(KEYINPUT59), .B(n588), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .Z(n593) );
  INV_X1 U655 ( .A(n591), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n596), .A2(n395), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U658 ( .A1(n596), .A2(n594), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U660 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n598) );
  NAND2_X1 U661 ( .A1(n596), .A2(n499), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

