//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1154, new_n1155,
    new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n450), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G113), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n472), .A2(new_n466), .A3(KEYINPUT69), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n472), .B2(new_n466), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n471), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n469), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NOR2_X1   g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n488), .B2(G112), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n487), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  OAI21_X1  g070(.A(G2104), .B1(new_n488), .B2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n463), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT71), .B1(new_n463), .B2(G2104), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n476), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT72), .B1(new_n469), .B2(new_n500), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n488), .A2(G138), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n469), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n469), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n508), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT74), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n523), .A2(G88), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G62), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n517), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G166));
  XOR2_X1   g112(.A(KEYINPUT76), .B(G89), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n530), .A2(new_n538), .B1(G63), .B2(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n517), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n529), .A2(new_n532), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n541), .B1(G51), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XOR2_X1   g119(.A(new_n544), .B(KEYINPUT7), .Z(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  NOR2_X1   g123(.A1(new_n529), .A2(new_n540), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n542), .A2(G52), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n518), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n540), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n542), .A2(G43), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n549), .A2(G81), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n542), .A2(G53), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n568), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n542), .A2(G53), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n540), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n549), .A2(G91), .B1(new_n576), .B2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n569), .A2(new_n578), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(G299));
  AND2_X1   g155(.A1(new_n535), .A2(new_n536), .ZN(G303));
  NAND2_X1  g156(.A1(new_n542), .A2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n549), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n542), .A2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n549), .A2(G86), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n517), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT79), .Z(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n549), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n542), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n518), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(new_n549), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n540), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n542), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT10), .B1(new_n604), .B2(new_n605), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT81), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n486), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n490), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n488), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n488), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n649), .B(new_n652), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT85), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(KEYINPUT17), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  INV_X1    g240(.A(new_n656), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n658), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n656), .A3(new_n658), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n632), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(G2100), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(G2100), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT89), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(new_n681), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n684), .A3(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n688), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT90), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  XNOR2_X1  g271(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G34), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n483), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G2084), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT98), .ZN(new_n704));
  OR2_X1    g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n486), .A2(G129), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n490), .A2(G141), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n488), .A2(G105), .A3(G2104), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND4_X1  g285(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n699), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G2072), .ZN(new_n715));
  OR2_X1    g290(.A1(G29), .A2(G33), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n490), .A2(G139), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n488), .A2(G103), .A3(G2104), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT25), .Z(new_n719));
  INV_X1    g294(.A(G127), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n478), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n717), .B(new_n719), .C1(new_n488), .C2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n699), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n714), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  NAND2_X1  g301(.A1(G171), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G5), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n704), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n699), .B1(new_n732), .B2(G28), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(G28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n738), .B1(new_n699), .B2(new_n631), .C1(new_n724), .C2(new_n715), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n701), .A2(new_n702), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n731), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G21), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G168), .B2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1966), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n699), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT99), .B(G2078), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n728), .A2(new_n729), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n741), .A2(new_n744), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n750), .A2(new_n731), .A3(new_n739), .A4(new_n740), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n755), .A2(KEYINPUT100), .A3(new_n744), .A4(new_n748), .ZN(new_n756));
  INV_X1    g331(.A(G16), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n757), .A2(KEYINPUT23), .A3(G20), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n759));
  INV_X1    g334(.A(G20), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(G16), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n761), .C1(new_n617), .C2(new_n757), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n699), .A2(G26), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n490), .A2(KEYINPUT94), .A3(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n486), .A2(G128), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n489), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n488), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n766), .A2(new_n767), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n765), .B1(new_n773), .B2(G29), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n765), .B(new_n774), .S(KEYINPUT28), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n754), .A2(new_n756), .A3(new_n764), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G22), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G166), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n757), .B1(new_n535), .B2(new_n536), .ZN(new_n782));
  OAI21_X1  g357(.A(G1971), .B1(new_n782), .B2(new_n778), .ZN(new_n783));
  MUX2_X1   g358(.A(G23), .B(G288), .S(G16), .Z(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(KEYINPUT33), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(KEYINPUT33), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n781), .A2(new_n783), .B1(new_n787), .B2(G1976), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n757), .B1(new_n594), .B2(new_n596), .ZN(new_n789));
  NOR2_X1   g364(.A1(G6), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT32), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n790), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n690), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1976), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n785), .B2(new_n786), .ZN(new_n796));
  INV_X1    g371(.A(new_n793), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n797), .A2(G1981), .A3(new_n791), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n788), .A2(new_n794), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT92), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G1986), .Z(new_n804));
  AND3_X1   g379(.A1(new_n799), .A2(KEYINPUT93), .A3(KEYINPUT34), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT93), .B1(new_n799), .B2(KEYINPUT34), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n801), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n486), .A2(G119), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n490), .A2(G131), .ZN(new_n809));
  NOR2_X1   g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(new_n488), .B2(G107), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT91), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT36), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n794), .A2(new_n798), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n781), .A2(new_n783), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n787), .A2(G1976), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(new_n821), .A3(new_n796), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n799), .A2(KEYINPUT93), .A3(KEYINPUT34), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n800), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  INV_X1    g403(.A(new_n816), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n804), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n777), .B1(new_n817), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n757), .A2(G19), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n561), .B2(new_n757), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1341), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n757), .A2(G4), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n613), .B2(new_n757), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1348), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n699), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n699), .ZN(new_n839));
  MUX2_X1   g414(.A(new_n838), .B(new_n839), .S(KEYINPUT101), .Z(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT29), .B(G2090), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n840), .B(new_n841), .Z(new_n842));
  NAND4_X1  g417(.A1(new_n831), .A2(new_n834), .A3(new_n837), .A4(new_n842), .ZN(G150));
  NAND2_X1  g418(.A1(G150), .A2(KEYINPUT102), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n845), .B(new_n777), .C1(new_n817), .C2(new_n830), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n834), .A4(new_n837), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n549), .A2(G93), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n542), .A2(G55), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n850), .B(new_n851), .C1(new_n518), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n612), .A2(new_n620), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT39), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n561), .B(new_n853), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n860), .B(new_n861), .Z(new_n862));
  OAI21_X1  g437(.A(new_n856), .B1(new_n862), .B2(G860), .ZN(G145));
  XNOR2_X1  g438(.A(new_n483), .B(new_n494), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  NOR2_X1   g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(new_n488), .B2(G118), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n489), .A2(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G130), .B2(new_n486), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n631), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n864), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n812), .B(new_n711), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n773), .B(new_n723), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n871), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n513), .A2(new_n515), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n503), .A2(new_n504), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n469), .A2(KEYINPUT72), .A3(new_n500), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT105), .B1(new_n879), .B2(new_n499), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n881), .B(new_n498), .C1(new_n877), .C2(new_n878), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n876), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n635), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n875), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT106), .B(G37), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT107), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n613), .ZN(new_n890));
  NAND2_X1  g465(.A1(G299), .A2(new_n612), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(KEYINPUT108), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n892), .B(KEYINPUT41), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(KEYINPUT108), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n623), .B(new_n861), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n893), .B2(new_n898), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(G166), .B(new_n597), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G288), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n903), .B(new_n904), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(new_n902), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n901), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n901), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G868), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n853), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n915), .ZN(G331));
  XNOR2_X1  g492(.A(new_n861), .B(G301), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G168), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n895), .C1(new_n896), .C2(KEYINPUT108), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n918), .B(G286), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n893), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n909), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  INV_X1    g500(.A(new_n909), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n926), .A3(new_n922), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n919), .A2(new_n896), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n919), .A2(new_n892), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n909), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n927), .A3(new_n886), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n928), .A2(new_n939), .A3(KEYINPUT43), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n933), .A2(new_n927), .A3(new_n929), .A4(new_n886), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n938), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n936), .B1(new_n944), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g520(.A(KEYINPUT53), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2078), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G164), .B2(G1384), .ZN(new_n951));
  OAI211_X1 g526(.A(G40), .B(new_n471), .C1(new_n481), .C2(new_n482), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n883), .A2(new_n955), .A3(new_n947), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n953), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n946), .A2(new_n954), .B1(new_n958), .B2(new_n729), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n498), .B1(new_n877), .B2(new_n878), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n876), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n883), .B2(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(G164), .A2(new_n950), .A3(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n952), .B1(new_n966), .B2(KEYINPUT116), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n946), .A2(G2078), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n959), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT122), .B1(new_n970), .B2(G171), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT122), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(G301), .C1(new_n959), .C2(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n507), .A2(new_n881), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n960), .A2(KEYINPUT105), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n977), .B2(new_n876), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n471), .B(new_n968), .C1(new_n978), .C2(KEYINPUT45), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n480), .A2(G40), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n948), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n974), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n948), .A2(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(new_n968), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n883), .A2(new_n947), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n950), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n983), .A2(KEYINPUT123), .A3(new_n986), .A4(new_n471), .ZN(new_n987));
  AND4_X1   g562(.A1(G301), .A2(new_n959), .A3(new_n982), .A4(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n971), .A2(new_n973), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT124), .B1(new_n989), .B2(KEYINPUT54), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT121), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT51), .ZN(new_n992));
  AOI21_X1  g567(.A(G1966), .B1(new_n965), .B2(new_n967), .ZN(new_n993));
  NOR2_X1   g568(.A1(KEYINPUT117), .A2(G2084), .ZN(new_n994));
  AND2_X1   g569(.A1(KEYINPUT117), .A2(G2084), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n958), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(G8), .B(new_n992), .C1(new_n997), .C2(G286), .ZN(new_n998));
  INV_X1    g573(.A(new_n992), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n991), .A2(KEYINPUT51), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n993), .A2(new_n996), .A3(G286), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(G8), .A3(G286), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n959), .A2(new_n982), .A3(new_n987), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G171), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n959), .A2(G301), .A3(new_n969), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(KEYINPUT54), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n948), .A2(new_n953), .A3(new_n951), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n1012), .B2(G1971), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1014), .A3(new_n780), .ZN(new_n1015));
  INV_X1    g590(.A(new_n958), .ZN(new_n1016));
  INV_X1    g591(.A(G2090), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(G8), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n985), .A2(new_n952), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n1002), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n795), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1025), .B(new_n1026), .C1(new_n795), .C2(G288), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n978), .A2(new_n953), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(new_n795), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n595), .B(new_n690), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1025), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1027), .A2(new_n1031), .A3(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1020), .B(KEYINPUT55), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n978), .A2(new_n955), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n961), .A2(new_n955), .A3(new_n947), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n953), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(new_n1017), .B1(new_n1011), .B2(new_n780), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n1044), .B2(new_n1002), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1023), .A2(new_n1038), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1010), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n970), .A2(G171), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n972), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n970), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n959), .A2(new_n982), .A3(new_n987), .A4(G301), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n990), .A2(new_n1005), .A3(new_n1047), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT125), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n577), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n577), .A2(new_n1060), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n572), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT119), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n763), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1012), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1059), .A2(new_n1070), .A3(new_n1064), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1069), .A2(new_n1067), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1066), .A2(new_n1076), .A3(new_n1071), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1016), .A2(G1348), .B1(G2067), .B2(new_n1028), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1080), .A2(new_n613), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1072), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n613), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT58), .B(G1341), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1011), .A2(G1996), .B1(new_n1024), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n561), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT59), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1078), .B2(new_n1072), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1072), .A2(new_n1089), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1075), .B2(new_n1073), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1084), .B(new_n1088), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1082), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1023), .A2(new_n1038), .A3(new_n1045), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1005), .A2(new_n1096), .A3(new_n1009), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT125), .A3(new_n990), .A4(new_n1055), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1058), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AND4_X1   g674(.A1(G8), .A2(new_n1038), .A3(new_n1022), .A4(new_n1019), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1037), .A2(new_n795), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(G288), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n592), .A2(new_n690), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1029), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1023), .A2(new_n1038), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n997), .A2(G8), .A3(G168), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1022), .B1(new_n1019), .B2(G8), .ZN(new_n1108));
  OR4_X1    g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1046), .B2(new_n1107), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1100), .B(new_n1104), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1046), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(KEYINPUT62), .B2(new_n1005), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT126), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1112), .B(new_n1116), .C1(KEYINPUT62), .C2(new_n1005), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1099), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n773), .B(G2067), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT112), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n711), .B(G1996), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n812), .A2(new_n815), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n812), .A2(new_n815), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n963), .A2(new_n953), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(G290), .B(G1986), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT113), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1119), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1126), .B(KEYINPUT127), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n773), .A2(G2067), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1128), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1129), .B1(new_n1122), .B2(new_n711), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1128), .B2(G1996), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n1128), .A2(new_n1140), .A3(G1996), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT47), .Z(new_n1144));
  NOR3_X1   g719(.A1(new_n1128), .A2(G1986), .A3(G290), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT48), .Z(new_n1146));
  AOI211_X1 g721(.A(new_n1138), .B(new_n1144), .C1(new_n1130), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1134), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g723(.A1(new_n887), .A2(G229), .ZN(new_n1150));
  INV_X1    g724(.A(new_n1150), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n672), .A2(new_n461), .A3(new_n654), .A4(new_n673), .ZN(new_n1152));
  NOR3_X1   g726(.A1(new_n944), .A2(new_n1151), .A3(new_n1152), .ZN(G308));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1154));
  AND2_X1   g728(.A1(new_n938), .A2(new_n940), .ZN(new_n1155));
  AND2_X1   g729(.A1(new_n942), .A2(new_n943), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n1150), .B(new_n1154), .C1(new_n1155), .C2(new_n1156), .ZN(G225));
endmodule


