

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759;

  XNOR2_X1 U368 ( .A(n428), .B(n358), .ZN(n658) );
  NOR2_X1 U369 ( .A1(n376), .A2(n694), .ZN(n455) );
  INV_X1 U370 ( .A(n681), .ZN(n609) );
  XNOR2_X1 U371 ( .A(n541), .B(KEYINPUT1), .ZN(n599) );
  NAND2_X2 U372 ( .A1(n368), .A2(n709), .ZN(n706) );
  NOR2_X1 U373 ( .A1(G902), .A2(n653), .ZN(n463) );
  XNOR2_X1 U374 ( .A(n743), .B(n440), .ZN(n462) );
  BUF_X2 U375 ( .A(n658), .Z(n391) );
  XNOR2_X2 U376 ( .A(n426), .B(n439), .ZN(n743) );
  XNOR2_X1 U377 ( .A(KEYINPUT3), .B(G113), .ZN(n447) );
  BUF_X1 U378 ( .A(G128), .Z(n390) );
  OR2_X1 U379 ( .A1(n646), .A2(n433), .ZN(n348) );
  NOR2_X1 U380 ( .A1(n658), .A2(n757), .ZN(n590) );
  NOR2_X1 U381 ( .A1(G953), .A2(G237), .ZN(n489) );
  XNOR2_X1 U382 ( .A(n447), .B(G101), .ZN(n350) );
  INV_X1 U383 ( .A(G146), .ZN(n440) );
  INV_X1 U384 ( .A(KEYINPUT22), .ZN(n387) );
  NAND2_X1 U385 ( .A1(n565), .A2(n564), .ZN(n396) );
  XNOR2_X1 U386 ( .A(n621), .B(n393), .ZN(n622) );
  XNOR2_X1 U387 ( .A(n589), .B(n588), .ZN(n637) );
  XNOR2_X1 U388 ( .A(n361), .B(KEYINPUT111), .ZN(n756) );
  AND2_X1 U389 ( .A1(n411), .A2(n352), .ZN(n410) );
  XNOR2_X1 U390 ( .A(n506), .B(n505), .ZN(n552) );
  XNOR2_X1 U391 ( .A(n665), .B(n373), .ZN(n646) );
  XNOR2_X1 U392 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U393 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U394 ( .A(n356), .ZN(n371) );
  XNOR2_X1 U395 ( .A(n525), .B(n524), .ZN(n665) );
  INV_X1 U396 ( .A(n350), .ZN(n518) );
  INV_X2 U397 ( .A(G953), .ZN(n745) );
  XNOR2_X1 U398 ( .A(n543), .B(KEYINPUT19), .ZN(n349) );
  XNOR2_X1 U399 ( .A(n543), .B(KEYINPUT19), .ZN(n384) );
  XNOR2_X2 U400 ( .A(n421), .B(n420), .ZN(n692) );
  NAND2_X1 U401 ( .A1(n379), .A2(n378), .ZN(n377) );
  AND2_X1 U402 ( .A1(n364), .A2(n360), .ZN(n378) );
  INV_X1 U403 ( .A(n756), .ZN(n360) );
  XNOR2_X1 U404 ( .A(G134), .B(G131), .ZN(n439) );
  NAND2_X1 U405 ( .A1(n538), .A2(n709), .ZN(n540) );
  AND2_X1 U406 ( .A1(n587), .A2(n354), .ZN(n538) );
  XNOR2_X1 U407 ( .A(G122), .B(G104), .ZN(n523) );
  NAND2_X1 U408 ( .A1(n419), .A2(n400), .ZN(n416) );
  NAND2_X1 U409 ( .A1(n385), .A2(n626), .ZN(n419) );
  NAND2_X1 U410 ( .A1(n699), .A2(n403), .ZN(n402) );
  INV_X1 U411 ( .A(KEYINPUT65), .ZN(n403) );
  INV_X1 U412 ( .A(G902), .ZN(n450) );
  XNOR2_X1 U413 ( .A(G137), .B(G119), .ZN(n444) );
  INV_X1 U414 ( .A(KEYINPUT68), .ZN(n443) );
  XOR2_X1 U415 ( .A(G116), .B(KEYINPUT5), .Z(n442) );
  AND2_X1 U416 ( .A1(n616), .A2(n394), .ZN(n620) );
  NOR2_X1 U417 ( .A1(n611), .A2(n610), .ZN(n616) );
  XNOR2_X1 U418 ( .A(n405), .B(G146), .ZN(n529) );
  INV_X1 U419 ( .A(G125), .ZN(n405) );
  XNOR2_X1 U420 ( .A(n561), .B(KEYINPUT38), .ZN(n549) );
  NAND2_X1 U421 ( .A1(n628), .A2(n434), .ZN(n433) );
  INV_X1 U422 ( .A(n533), .ZN(n434) );
  INV_X1 U423 ( .A(KEYINPUT108), .ZN(n407) );
  XNOR2_X1 U424 ( .A(n353), .B(n476), .ZN(n587) );
  XNOR2_X1 U425 ( .A(n377), .B(n359), .ZN(n565) );
  XNOR2_X1 U426 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n492) );
  XNOR2_X1 U427 ( .A(G113), .B(G143), .ZN(n498) );
  XNOR2_X1 U428 ( .A(n529), .B(n404), .ZN(n490) );
  INV_X1 U429 ( .A(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U430 ( .A(n431), .B(n430), .ZN(n386) );
  XNOR2_X1 U431 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U432 ( .A1(n586), .A2(KEYINPUT102), .ZN(n413) );
  XNOR2_X1 U433 ( .A(n536), .B(KEYINPUT100), .ZN(n537) );
  INV_X1 U434 ( .A(KEYINPUT6), .ZN(n536) );
  INV_X1 U435 ( .A(n587), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U437 ( .A(n458), .B(n436), .ZN(n460) );
  INV_X1 U438 ( .A(G469), .ZN(n418) );
  AND2_X1 U439 ( .A1(n633), .A2(G953), .ZN(n742) );
  INV_X1 U440 ( .A(n709), .ZN(n367) );
  INV_X1 U441 ( .A(KEYINPUT46), .ZN(n380) );
  AND2_X1 U442 ( .A1(n544), .A2(n365), .ZN(n364) );
  XNOR2_X1 U443 ( .A(n401), .B(KEYINPUT47), .ZN(n365) );
  NOR2_X1 U444 ( .A1(n679), .A2(n402), .ZN(n401) );
  NOR2_X1 U445 ( .A1(n676), .A2(n670), .ZN(n394) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n479) );
  AND2_X1 U447 ( .A1(n613), .A2(n566), .ZN(n567) );
  INV_X1 U448 ( .A(n694), .ZN(n372) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n557) );
  INV_X1 U450 ( .A(KEYINPUT80), .ZN(n393) );
  XNOR2_X1 U451 ( .A(G131), .B(KEYINPUT96), .ZN(n494) );
  NOR2_X1 U452 ( .A1(n659), .A2(n628), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n396), .B(KEYINPUT69), .ZN(n366) );
  INV_X1 U454 ( .A(G237), .ZN(n437) );
  INV_X1 U455 ( .A(KEYINPUT88), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n462), .B(n449), .ZN(n630) );
  XNOR2_X1 U457 ( .A(n522), .B(n369), .ZN(n467) );
  INV_X1 U458 ( .A(n390), .ZN(n369) );
  XOR2_X1 U459 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n466) );
  XOR2_X1 U460 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n508) );
  XNOR2_X1 U461 ( .A(G134), .B(G122), .ZN(n507) );
  XNOR2_X1 U462 ( .A(G101), .B(G104), .ZN(n456) );
  XOR2_X1 U463 ( .A(G110), .B(KEYINPUT83), .Z(n457) );
  XOR2_X1 U464 ( .A(G107), .B(KEYINPUT89), .Z(n436) );
  XNOR2_X1 U465 ( .A(G137), .B(G140), .ZN(n470) );
  INV_X1 U466 ( .A(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U467 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n527) );
  INV_X1 U468 ( .A(KEYINPUT70), .ZN(n420) );
  NOR2_X1 U469 ( .A1(n539), .A2(n540), .ZN(n558) );
  NAND2_X1 U470 ( .A1(n348), .A2(n351), .ZN(n561) );
  AND2_X1 U471 ( .A1(n488), .A2(n487), .ZN(n545) );
  XNOR2_X1 U472 ( .A(KEYINPUT106), .B(n453), .ZN(n454) );
  XNOR2_X1 U473 ( .A(n408), .B(n406), .ZN(n542) );
  XNOR2_X1 U474 ( .A(n407), .B(KEYINPUT28), .ZN(n406) );
  XOR2_X1 U475 ( .A(n630), .B(KEYINPUT62), .Z(n631) );
  XNOR2_X1 U476 ( .A(n350), .B(n521), .ZN(n525) );
  XNOR2_X1 U477 ( .A(n502), .B(n501), .ZN(n639) );
  XNOR2_X1 U478 ( .A(n548), .B(KEYINPUT40), .ZN(n758) );
  NAND2_X1 U479 ( .A1(n362), .A2(n586), .ZN(n361) );
  XNOR2_X1 U480 ( .A(n422), .B(n363), .ZN(n362) );
  INV_X1 U481 ( .A(KEYINPUT36), .ZN(n363) );
  NAND2_X1 U482 ( .A1(n386), .A2(n429), .ZN(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT32), .B(n585), .ZN(n757) );
  NAND2_X1 U484 ( .A1(n410), .A2(n409), .ZN(n589) );
  NAND2_X1 U485 ( .A1(n414), .A2(n413), .ZN(n409) );
  NAND2_X1 U486 ( .A1(n609), .A2(n618), .ZN(n671) );
  NOR2_X1 U487 ( .A1(n656), .A2(n742), .ZN(n657) );
  NOR2_X1 U488 ( .A1(n389), .A2(n356), .ZN(n351) );
  AND2_X1 U489 ( .A1(n412), .A2(n357), .ZN(n352) );
  XNOR2_X1 U490 ( .A(KEYINPUT15), .B(G902), .ZN(n628) );
  XOR2_X1 U491 ( .A(n475), .B(KEYINPUT90), .Z(n353) );
  XOR2_X1 U492 ( .A(KEYINPUT74), .B(n486), .Z(n354) );
  XNOR2_X1 U493 ( .A(n438), .B(KEYINPUT85), .ZN(n694) );
  NOR2_X1 U494 ( .A1(n395), .A2(n606), .ZN(n355) );
  AND2_X1 U495 ( .A1(n629), .A2(n533), .ZN(n356) );
  AND2_X1 U496 ( .A1(n376), .A2(n587), .ZN(n357) );
  XOR2_X1 U497 ( .A(n580), .B(KEYINPUT72), .Z(n358) );
  XNOR2_X1 U498 ( .A(n557), .B(KEYINPUT78), .ZN(n359) );
  INV_X1 U499 ( .A(n628), .ZN(n629) );
  NAND2_X1 U500 ( .A1(n382), .A2(n366), .ZN(n385) );
  NAND2_X1 U501 ( .A1(n627), .A2(n366), .ZN(n397) );
  AND2_X1 U502 ( .A1(n587), .A2(n367), .ZN(n711) );
  NOR2_X1 U503 ( .A1(n581), .A2(n368), .ZN(n582) );
  NAND2_X1 U504 ( .A1(n707), .A2(n368), .ZN(n612) );
  XNOR2_X2 U505 ( .A(G119), .B(G110), .ZN(n522) );
  AND2_X2 U506 ( .A1(n646), .A2(n533), .ZN(n389) );
  XNOR2_X1 U507 ( .A(n712), .B(n537), .ZN(n613) );
  XNOR2_X1 U508 ( .A(n712), .B(KEYINPUT101), .ZN(n376) );
  BUF_X1 U509 ( .A(n712), .Z(n395) );
  NOR2_X1 U510 ( .A1(n389), .A2(n370), .ZN(n432) );
  XNOR2_X1 U511 ( .A(n530), .B(n531), .ZN(n373) );
  NOR2_X2 U512 ( .A1(n374), .A2(n583), .ZN(n388) );
  NOR2_X1 U513 ( .A1(n717), .A2(n374), .ZN(n601) );
  XNOR2_X1 U514 ( .A(n374), .B(n392), .ZN(n383) );
  XNOR2_X2 U515 ( .A(n578), .B(n577), .ZN(n374) );
  XNOR2_X2 U516 ( .A(n375), .B(n569), .ZN(n704) );
  NAND2_X1 U517 ( .A1(n567), .A2(n568), .ZN(n375) );
  NOR2_X1 U518 ( .A1(n540), .A2(n376), .ZN(n408) );
  XNOR2_X1 U519 ( .A(n381), .B(n380), .ZN(n379) );
  NAND2_X1 U520 ( .A1(n758), .A2(n759), .ZN(n381) );
  NAND2_X1 U521 ( .A1(n704), .A2(n383), .ZN(n431) );
  NAND2_X1 U522 ( .A1(n355), .A2(n383), .ZN(n608) );
  NAND2_X1 U523 ( .A1(n384), .A2(n575), .ZN(n578) );
  NAND2_X1 U524 ( .A1(n554), .A2(n349), .ZN(n679) );
  AND2_X2 U525 ( .A1(n415), .A2(n416), .ZN(n738) );
  XNOR2_X2 U526 ( .A(n388), .B(n387), .ZN(n614) );
  NAND2_X1 U527 ( .A1(n738), .A2(G210), .ZN(n648) );
  INV_X1 U528 ( .A(n579), .ZN(n429) );
  NAND2_X1 U529 ( .A1(n738), .A2(G475), .ZN(n641) );
  NAND2_X2 U530 ( .A1(n432), .A2(n348), .ZN(n543) );
  NOR2_X2 U531 ( .A1(n634), .A2(n742), .ZN(n636) );
  NOR2_X2 U532 ( .A1(n642), .A2(n742), .ZN(n643) );
  NOR2_X2 U533 ( .A1(n649), .A2(n742), .ZN(n650) );
  XNOR2_X2 U534 ( .A(n452), .B(n451), .ZN(n712) );
  NOR2_X2 U535 ( .A1(n659), .A2(n396), .ZN(n689) );
  INV_X1 U536 ( .A(n692), .ZN(n415) );
  XNOR2_X1 U537 ( .A(n396), .B(n747), .ZN(n746) );
  NAND2_X1 U538 ( .A1(n397), .A2(n399), .ZN(n398) );
  NAND2_X1 U539 ( .A1(n398), .A2(n629), .ZN(n400) );
  INV_X1 U540 ( .A(KEYINPUT2), .ZN(n399) );
  NAND2_X1 U541 ( .A1(n614), .A2(KEYINPUT102), .ZN(n411) );
  NAND2_X1 U542 ( .A1(n586), .A2(KEYINPUT102), .ZN(n412) );
  INV_X1 U543 ( .A(n614), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n689), .A2(KEYINPUT2), .ZN(n421) );
  NAND2_X1 U545 ( .A1(n417), .A2(n416), .ZN(n655) );
  NOR2_X1 U546 ( .A1(n692), .A2(n418), .ZN(n417) );
  XNOR2_X2 U547 ( .A(n512), .B(n427), .ZN(n426) );
  NAND2_X1 U548 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U549 ( .A(n543), .ZN(n423) );
  XNOR2_X1 U550 ( .A(n558), .B(KEYINPUT110), .ZN(n424) );
  XNOR2_X1 U551 ( .A(n426), .B(n425), .ZN(n530) );
  INV_X1 U552 ( .A(n529), .ZN(n425) );
  INV_X1 U553 ( .A(KEYINPUT34), .ZN(n430) );
  XNOR2_X2 U554 ( .A(G116), .B(G107), .ZN(n520) );
  XNOR2_X1 U555 ( .A(n462), .B(n461), .ZN(n653) );
  AND2_X1 U556 ( .A1(G227), .A2(n745), .ZN(n435) );
  INV_X1 U557 ( .A(KEYINPUT76), .ZN(n626) );
  XNOR2_X1 U558 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U559 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U560 ( .A(n435), .B(n470), .ZN(n459) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  AND2_X1 U562 ( .A1(n605), .A2(n354), .ZN(n487) );
  NAND2_X1 U563 ( .A1(n450), .A2(n437), .ZN(n532) );
  NAND2_X1 U564 ( .A1(n532), .A2(G214), .ZN(n438) );
  XNOR2_X2 U565 ( .A(G143), .B(G128), .ZN(n512) );
  NAND2_X1 U566 ( .A1(n489), .A2(G210), .ZN(n441) );
  XNOR2_X1 U567 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U568 ( .A(n518), .B(n448), .ZN(n449) );
  NAND2_X1 U569 ( .A1(n630), .A2(n450), .ZN(n452) );
  XOR2_X1 U570 ( .A(G472), .B(KEYINPUT91), .Z(n451) );
  XOR2_X1 U571 ( .A(KEYINPUT105), .B(KEYINPUT30), .Z(n453) );
  XNOR2_X1 U572 ( .A(n455), .B(n454), .ZN(n488) );
  XNOR2_X1 U573 ( .A(KEYINPUT66), .B(G469), .ZN(n464) );
  XNOR2_X1 U574 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X2 U575 ( .A(n464), .B(n463), .ZN(n541) );
  NAND2_X1 U576 ( .A1(G234), .A2(n745), .ZN(n465) );
  XOR2_X1 U577 ( .A(KEYINPUT8), .B(n465), .Z(n509) );
  NAND2_X1 U578 ( .A1(n509), .A2(G221), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U580 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U581 ( .A(n490), .B(n470), .ZN(n744) );
  XNOR2_X1 U582 ( .A(n471), .B(n744), .ZN(n739) );
  NOR2_X1 U583 ( .A1(n739), .A2(G902), .ZN(n476) );
  XOR2_X1 U584 ( .A(KEYINPUT25), .B(KEYINPUT71), .Z(n474) );
  NAND2_X1 U585 ( .A1(n628), .A2(G234), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n472), .B(KEYINPUT20), .ZN(n477) );
  NAND2_X1 U587 ( .A1(n477), .A2(G217), .ZN(n473) );
  XNOR2_X1 U588 ( .A(n474), .B(n473), .ZN(n475) );
  AND2_X1 U589 ( .A1(n477), .A2(G221), .ZN(n478) );
  XNOR2_X1 U590 ( .A(n478), .B(KEYINPUT21), .ZN(n709) );
  NOR2_X1 U591 ( .A1(n541), .A2(n706), .ZN(n605) );
  XNOR2_X1 U592 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U593 ( .A1(G952), .A2(n481), .ZN(n480) );
  XOR2_X1 U594 ( .A(KEYINPUT86), .B(n480), .Z(n724) );
  NAND2_X1 U595 ( .A1(n745), .A2(n724), .ZN(n573) );
  INV_X1 U596 ( .A(n573), .ZN(n485) );
  NAND2_X1 U597 ( .A1(G902), .A2(n481), .ZN(n570) );
  NOR2_X1 U598 ( .A1(G900), .A2(n570), .ZN(n482) );
  NAND2_X1 U599 ( .A1(G953), .A2(n482), .ZN(n483) );
  XOR2_X1 U600 ( .A(KEYINPUT104), .B(n483), .Z(n484) );
  NOR2_X1 U601 ( .A1(n485), .A2(n484), .ZN(n486) );
  NAND2_X1 U602 ( .A1(G214), .A2(n489), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n491), .B(n490), .ZN(n502) );
  XOR2_X1 U604 ( .A(KEYINPUT95), .B(G140), .Z(n493) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U606 ( .A(KEYINPUT97), .B(KEYINPUT94), .Z(n495) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n497), .B(n496), .ZN(n500) );
  XOR2_X1 U609 ( .A(n498), .B(n523), .Z(n499) );
  NOR2_X1 U610 ( .A1(G902), .A2(n639), .ZN(n506) );
  XNOR2_X1 U611 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n504) );
  INV_X1 U612 ( .A(G475), .ZN(n503) );
  INV_X1 U613 ( .A(n552), .ZN(n517) );
  XNOR2_X1 U614 ( .A(KEYINPUT99), .B(G478), .ZN(n516) );
  XNOR2_X1 U615 ( .A(n508), .B(n507), .ZN(n511) );
  NAND2_X1 U616 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n511), .B(n510), .ZN(n514) );
  XOR2_X1 U618 ( .A(n512), .B(n520), .Z(n513) );
  XNOR2_X1 U619 ( .A(n514), .B(n513), .ZN(n735) );
  NOR2_X1 U620 ( .A1(G902), .A2(n735), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n550) );
  NAND2_X1 U622 ( .A1(n517), .A2(n550), .ZN(n579) );
  XNOR2_X1 U623 ( .A(KEYINPUT83), .B(KEYINPUT16), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n745), .A2(G224), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n526), .B(KEYINPUT84), .ZN(n528) );
  XNOR2_X1 U628 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n532), .A2(G210), .ZN(n533) );
  NOR2_X1 U630 ( .A1(n579), .A2(n561), .ZN(n534) );
  NAND2_X1 U631 ( .A1(n545), .A2(n534), .ZN(n535) );
  XNOR2_X1 U632 ( .A(KEYINPUT107), .B(n535), .ZN(n752) );
  XNOR2_X1 U633 ( .A(n752), .B(KEYINPUT75), .ZN(n544) );
  OR2_X1 U634 ( .A1(n552), .A2(n550), .ZN(n681) );
  NAND2_X1 U635 ( .A1(n609), .A2(n613), .ZN(n539) );
  INV_X1 U636 ( .A(n599), .ZN(n586) );
  INV_X1 U637 ( .A(n586), .ZN(n707) );
  NOR2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n554) );
  NAND2_X1 U639 ( .A1(n552), .A2(n550), .ZN(n684) );
  NAND2_X1 U640 ( .A1(n684), .A2(n681), .ZN(n699) );
  NAND2_X1 U641 ( .A1(n545), .A2(n549), .ZN(n547) );
  XOR2_X1 U642 ( .A(KEYINPUT79), .B(KEYINPUT39), .Z(n546) );
  XNOR2_X1 U643 ( .A(n547), .B(n546), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n563), .A2(n609), .ZN(n548) );
  XOR2_X1 U645 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n556) );
  INV_X1 U646 ( .A(n549), .ZN(n695) );
  NOR2_X1 U647 ( .A1(n695), .A2(n694), .ZN(n700) );
  INV_X1 U648 ( .A(n550), .ZN(n551) );
  AND2_X1 U649 ( .A1(n552), .A2(n551), .ZN(n697) );
  NAND2_X1 U650 ( .A1(n700), .A2(n697), .ZN(n553) );
  XNOR2_X1 U651 ( .A(n553), .B(KEYINPUT41), .ZN(n720) );
  NAND2_X1 U652 ( .A1(n720), .A2(n554), .ZN(n555) );
  XNOR2_X1 U653 ( .A(n556), .B(n555), .ZN(n759) );
  NAND2_X1 U654 ( .A1(n558), .A2(n707), .ZN(n559) );
  NOR2_X1 U655 ( .A1(n694), .A2(n559), .ZN(n560) );
  XOR2_X1 U656 ( .A(n560), .B(KEYINPUT43), .Z(n562) );
  NAND2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n687) );
  INV_X1 U658 ( .A(n684), .ZN(n617) );
  NAND2_X1 U659 ( .A1(n563), .A2(n617), .ZN(n686) );
  AND2_X1 U660 ( .A1(n687), .A2(n686), .ZN(n564) );
  INV_X1 U661 ( .A(n599), .ZN(n568) );
  INV_X1 U662 ( .A(n706), .ZN(n566) );
  XNOR2_X1 U663 ( .A(KEYINPUT82), .B(KEYINPUT33), .ZN(n569) );
  NOR2_X1 U664 ( .A1(G898), .A2(n745), .ZN(n666) );
  INV_X1 U665 ( .A(n570), .ZN(n571) );
  NAND2_X1 U666 ( .A1(n666), .A2(n571), .ZN(n572) );
  AND2_X1 U667 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n574), .B(KEYINPUT87), .ZN(n575) );
  INV_X1 U669 ( .A(KEYINPUT81), .ZN(n576) );
  XNOR2_X1 U670 ( .A(n576), .B(KEYINPUT0), .ZN(n577) );
  XNOR2_X1 U671 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n580) );
  OR2_X1 U672 ( .A1(n613), .A2(n599), .ZN(n581) );
  XNOR2_X1 U673 ( .A(n582), .B(KEYINPUT73), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n697), .A2(n709), .ZN(n583) );
  NOR2_X1 U675 ( .A1(n584), .A2(n614), .ZN(n585) );
  INV_X1 U676 ( .A(KEYINPUT103), .ZN(n588) );
  NAND2_X1 U677 ( .A1(n590), .A2(n637), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(n594), .ZN(n593) );
  INV_X1 U679 ( .A(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n598) );
  INV_X1 U681 ( .A(KEYINPUT67), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n594), .A2(KEYINPUT44), .ZN(n595) );
  NOR2_X1 U683 ( .A1(n757), .A2(n595), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n596), .A2(n637), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n623) );
  INV_X1 U686 ( .A(n699), .ZN(n604) );
  INV_X1 U687 ( .A(KEYINPUT31), .ZN(n602) );
  NOR2_X1 U688 ( .A1(n599), .A2(n706), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n395), .A2(n600), .ZN(n717) );
  XNOR2_X1 U690 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U691 ( .A(KEYINPUT93), .B(n603), .ZN(n683) );
  NOR2_X1 U692 ( .A1(n604), .A2(n683), .ZN(n611) );
  INV_X1 U693 ( .A(n605), .ZN(n606) );
  INV_X1 U694 ( .A(KEYINPUT92), .ZN(n607) );
  XNOR2_X1 U695 ( .A(n608), .B(n607), .ZN(n618) );
  INV_X1 U696 ( .A(n671), .ZN(n610) );
  OR2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n670) );
  AND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n676) );
  NAND2_X1 U700 ( .A1(n391), .A2(KEYINPUT44), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n624) );
  XNOR2_X2 U704 ( .A(n625), .B(n624), .ZN(n659) );
  NOR2_X1 U705 ( .A1(n659), .A2(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n738), .A2(G472), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U708 ( .A(G952), .ZN(n633) );
  INV_X1 U709 ( .A(KEYINPUT63), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(G57) );
  XNOR2_X1 U711 ( .A(n637), .B(G110), .ZN(G12) );
  XNOR2_X1 U712 ( .A(KEYINPUT127), .B(KEYINPUT59), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U715 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n644) );
  XOR2_X1 U716 ( .A(n644), .B(KEYINPUT55), .Z(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U720 ( .A(KEYINPUT125), .B(KEYINPUT57), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(KEYINPUT58), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(KEYINPUT126), .ZN(G54) );
  XOR2_X1 U725 ( .A(n391), .B(G122), .Z(G24) );
  INV_X1 U726 ( .A(n659), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n660), .A2(n745), .ZN(n664) );
  NAND2_X1 U728 ( .A1(G953), .A2(G224), .ZN(n661) );
  XNOR2_X1 U729 ( .A(KEYINPUT61), .B(n661), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n662), .A2(G898), .ZN(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n669) );
  INV_X1 U732 ( .A(n665), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n669), .B(n668), .ZN(G69) );
  XOR2_X1 U735 ( .A(G101), .B(n670), .Z(G3) );
  XNOR2_X1 U736 ( .A(G104), .B(KEYINPUT112), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(n671), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n674) );
  XNOR2_X1 U739 ( .A(G107), .B(KEYINPUT26), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n676), .B(n675), .ZN(G9) );
  NOR2_X1 U742 ( .A1(n679), .A2(n684), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n390), .B(KEYINPUT29), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n678), .B(n677), .ZN(G30) );
  NOR2_X1 U745 ( .A1(n679), .A2(n681), .ZN(n680) );
  XOR2_X1 U746 ( .A(G146), .B(n680), .Z(G48) );
  NOR2_X1 U747 ( .A1(n681), .A2(n683), .ZN(n682) );
  XOR2_X1 U748 ( .A(G113), .B(n682), .Z(G15) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U750 ( .A(G116), .B(n685), .Z(G18) );
  XNOR2_X1 U751 ( .A(G134), .B(n686), .ZN(G36) );
  XNOR2_X1 U752 ( .A(n687), .B(G140), .ZN(n688) );
  XNOR2_X1 U753 ( .A(KEYINPUT116), .B(n688), .ZN(G42) );
  XOR2_X1 U754 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n734) );
  BUF_X1 U755 ( .A(n689), .Z(n690) );
  NOR2_X1 U756 ( .A1(n690), .A2(KEYINPUT2), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n731) );
  NAND2_X1 U758 ( .A1(n720), .A2(n704), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT120), .ZN(n727) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U762 ( .A(n698), .B(KEYINPUT118), .ZN(n702) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U766 ( .A(KEYINPUT119), .B(n705), .Z(n722) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(KEYINPUT50), .B(n708), .ZN(n715) );
  XNOR2_X1 U769 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n713), .A2(n395), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT51), .B(n718), .Z(n719) );
  NAND2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT52), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT121), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(n745), .ZN(n730) );
  NOR2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n732), .B(KEYINPUT122), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(G75) );
  NAND2_X1 U785 ( .A1(n738), .A2(G478), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U787 ( .A1(n742), .A2(n737), .ZN(G63) );
  NAND2_X1 U788 ( .A1(n738), .A2(G217), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n742), .A2(n741), .ZN(G66) );
  XNOR2_X1 U791 ( .A(n743), .B(n744), .ZN(n747) );
  NAND2_X1 U792 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U793 ( .A(G227), .B(n747), .ZN(n748) );
  NAND2_X1 U794 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U795 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U796 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U797 ( .A(G143), .B(n752), .Z(G45) );
  XOR2_X1 U798 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n754) );
  XNOR2_X1 U799 ( .A(G125), .B(KEYINPUT115), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U801 ( .A(n756), .B(n755), .ZN(G27) );
  XOR2_X1 U802 ( .A(G119), .B(n757), .Z(G21) );
  XNOR2_X1 U803 ( .A(n758), .B(G131), .ZN(G33) );
  XNOR2_X1 U804 ( .A(G137), .B(n759), .ZN(G39) );
endmodule

