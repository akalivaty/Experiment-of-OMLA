//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(new_n189), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(G128), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n200), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n201), .B(G146), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n205), .B2(new_n209), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n199), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT11), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  OR3_X1    g033(.A1(new_n216), .A2(KEYINPUT66), .A3(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n216), .B2(G134), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n216), .A2(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n213), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n203), .A2(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n201), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n236), .A2(new_n238), .B1(new_n194), .B2(new_n232), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n218), .A2(new_n221), .A3(new_n220), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n222), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n197), .A2(new_n198), .B1(G143), .B2(new_n203), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT68), .B(new_n231), .C1(new_n245), .C2(new_n200), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n226), .B1(new_n248), .B2(new_n199), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n194), .A2(new_n232), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n231), .A2(new_n234), .A3(new_n237), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n237), .B1(new_n231), .B2(new_n234), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n253), .A2(KEYINPUT65), .B1(new_n222), .B2(new_n241), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n239), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n249), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n193), .B(new_n244), .C1(new_n257), .C2(KEYINPUT30), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n228), .A2(new_n192), .A3(new_n243), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n212), .A2(new_n227), .B1(new_n239), .B2(new_n242), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n192), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n254), .A2(new_n256), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n193), .B1(new_n274), .B2(new_n249), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n265), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n267), .A2(new_n268), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n270), .A2(new_n192), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n269), .B2(new_n272), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n266), .A2(new_n268), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n187), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n187), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n266), .B1(new_n270), .B2(new_n192), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n258), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n258), .A2(new_n289), .A3(new_n285), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n265), .B1(new_n273), .B2(new_n275), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n258), .B2(new_n285), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n284), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n282), .B1(KEYINPUT32), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  AOI211_X1 g112(.A(new_n292), .B(new_n294), .C1(new_n288), .C2(new_n290), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT71), .B(new_n298), .C1(new_n299), .C2(new_n284), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n297), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT16), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(G140), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT16), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n309), .A2(G146), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G125), .B(G140), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n203), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n200), .A2(KEYINPUT73), .A3(G119), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n319), .C1(G119), .C2(new_n200), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT74), .B1(new_n317), .B2(G128), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n324), .A2(KEYINPUT23), .B1(new_n317), .B2(G128), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(KEYINPUT23), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n326), .B2(G110), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n315), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n309), .A2(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n203), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n309), .A2(new_n312), .A3(G146), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n330), .B(new_n334), .C1(new_n322), .C2(new_n320), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n329), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n329), .B2(new_n335), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n340), .A2(new_n341), .A3(G902), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n304), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n341), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n329), .A2(new_n335), .A3(new_n339), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n283), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT72), .B(G217), .Z(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n283), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(G902), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n303), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  OAI21_X1  g170(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G104), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G104), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G107), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT80), .B(G101), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(G104), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT78), .B1(new_n367), .B2(KEYINPUT3), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n363), .C2(G107), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n365), .B(new_n366), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n364), .B2(new_n361), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(KEYINPUT10), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n199), .A2(new_n205), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n371), .A3(new_n372), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n373), .A2(new_n212), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n241), .A2(new_n222), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT3), .B1(new_n363), .B2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n369), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(KEYINPUT79), .A3(new_n365), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT79), .B1(new_n384), .B2(new_n365), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n380), .B1(new_n387), .B2(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n365), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(KEYINPUT79), .A3(new_n365), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n239), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n378), .B(new_n379), .C1(new_n388), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n337), .A2(G227), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n199), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n246), .B2(new_n247), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n371), .A2(new_n372), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n376), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT12), .B1(new_n406), .B2(new_n242), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n379), .C1(new_n405), .C2(new_n376), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n397), .B(new_n401), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n378), .B1(new_n388), .B2(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n242), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n401), .B1(new_n413), .B2(new_n397), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n359), .B(new_n283), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n397), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n385), .A2(new_n386), .A3(new_n393), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n239), .B(new_n395), .C1(new_n419), .C2(new_n380), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n379), .B1(new_n420), .B2(new_n378), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n400), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n422), .B2(new_n410), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n359), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n397), .B1(new_n407), .B2(new_n409), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n400), .B(KEYINPUT77), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n413), .A2(new_n397), .A3(new_n401), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n359), .B1(new_n430), .B2(new_n283), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n358), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n317), .A2(G116), .ZN(new_n436));
  OAI21_X1  g250(.A(G113), .B1(new_n436), .B2(KEYINPUT5), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n190), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n371), .A3(new_n372), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n395), .A2(new_n193), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n388), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n440), .B(new_n443), .C1(new_n388), .C2(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n403), .A2(new_n307), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n253), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n337), .A2(G224), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT82), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n452), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n452), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n454), .A2(new_n457), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n439), .A2(new_n404), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n443), .B(KEYINPUT8), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n437), .A2(KEYINPUT83), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n190), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n461), .B(new_n462), .C1(new_n465), .C2(new_n404), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n458), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n467), .B2(new_n446), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n456), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n456), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n434), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n456), .A2(new_n468), .ZN(new_n474));
  INV_X1    g288(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n456), .A2(new_n468), .A3(new_n469), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n434), .ZN(new_n480));
  NOR3_X1   g294(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n481));
  INV_X1    g295(.A(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G113), .ZN(new_n483));
  INV_X1    g297(.A(G113), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G122), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n485), .A3(G104), .ZN(new_n486));
  AOI21_X1  g300(.A(G104), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT19), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n305), .A2(G125), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n310), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT19), .ZN(new_n493));
  AOI21_X1  g307(.A(G146), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n489), .B1(new_n494), .B2(new_n313), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n261), .A2(G214), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n201), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n219), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G237), .ZN(new_n500));
  AND4_X1   g314(.A1(G143), .A2(new_n500), .A3(new_n337), .A4(G214), .ZN(new_n501));
  AOI21_X1  g315(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT19), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT19), .B1(new_n306), .B2(new_n308), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n203), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n333), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n314), .B(new_n203), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT18), .B(G131), .C1(new_n501), .C2(new_n502), .ZN(new_n511));
  NAND2_X1  g325(.A1(KEYINPUT18), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n497), .A2(new_n498), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n488), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT86), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n484), .A2(G122), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n482), .A2(G113), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n363), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n483), .A2(new_n485), .A3(G104), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n499), .A2(new_n503), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT17), .B(G131), .C1(new_n501), .C2(new_n502), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n332), .A2(new_n333), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n514), .B(new_n523), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n481), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT88), .B(new_n481), .C1(new_n515), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n535));
  OR3_X1    g349(.A1(new_n515), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n515), .B2(new_n529), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n534), .B1(KEYINPUT20), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G475), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n525), .A2(new_n527), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n528), .B1(new_n543), .B2(new_n488), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n283), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n349), .A2(G953), .A3(new_n356), .ZN(new_n546));
  XNOR2_X1  g360(.A(G116), .B(G122), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(new_n360), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n201), .A2(G128), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT13), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n200), .A2(G143), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(new_n550), .ZN(new_n554));
  OAI21_X1  g368(.A(G134), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(new_n552), .A3(new_n213), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G116), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT14), .A3(G122), .ZN(new_n559));
  INV_X1    g373(.A(new_n547), .ZN(new_n560));
  OAI211_X1 g374(.A(G107), .B(new_n559), .C1(new_n560), .C2(KEYINPUT14), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n549), .A2(new_n552), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G134), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n556), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n547), .A2(new_n360), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n546), .B1(new_n557), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n557), .A2(new_n566), .A3(new_n546), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n567), .B1(new_n572), .B2(KEYINPUT89), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n573), .A3(new_n283), .ZN(new_n574));
  INV_X1    g388(.A(G478), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n337), .A2(G952), .ZN(new_n578));
  INV_X1    g392(.A(G234), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n500), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n283), .B(new_n337), .C1(G234), .C2(G237), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n576), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n571), .A2(new_n573), .A3(new_n283), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n540), .A2(new_n545), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n433), .A2(new_n473), .A3(new_n480), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n355), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT90), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n366), .ZN(G3));
  NAND2_X1  g407(.A1(new_n291), .A2(new_n295), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n187), .B1(new_n594), .B2(new_n283), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n296), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n539), .A2(KEYINPUT20), .ZN(new_n597));
  INV_X1    g411(.A(new_n534), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n545), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n575), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n572), .B1(new_n603), .B2(new_n567), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n568), .A2(KEYINPUT91), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT33), .B1(new_n571), .B2(new_n573), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n574), .A2(new_n575), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n433), .A2(new_n596), .A3(new_n354), .A4(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n434), .B(new_n585), .C1(new_n470), .C2(new_n471), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  AND2_X1   g431(.A1(new_n536), .A2(new_n538), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n481), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n597), .ZN(new_n620));
  INV_X1    g434(.A(new_n545), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n577), .A2(new_n587), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(new_n354), .A3(new_n433), .A4(new_n596), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n360), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(new_n596), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n329), .A2(new_n335), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(KEYINPUT93), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(KEYINPUT93), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n339), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(KEYINPUT36), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI22_X1  g450(.A1(new_n632), .A2(new_n631), .B1(KEYINPUT36), .B2(new_n634), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n352), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n351), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n590), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT37), .B(G110), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT94), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n351), .A2(new_n638), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n434), .B(new_n644), .C1(new_n470), .C2(new_n471), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n581), .B1(new_n582), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n303), .A2(new_n433), .A3(new_n646), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(KEYINPUT95), .B(KEYINPUT39), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n648), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n433), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n656), .B(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n258), .A2(new_n285), .ZN(new_n663));
  INV_X1    g477(.A(new_n278), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n259), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n665), .B2(new_n265), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n187), .B1(new_n666), .B2(new_n283), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n300), .A2(new_n302), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n470), .A2(new_n471), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n600), .A2(new_n434), .A3(new_n622), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n670), .A2(new_n674), .A3(new_n644), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n660), .A2(new_n662), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  AOI21_X1  g492(.A(new_n431), .B1(new_n417), .B2(new_n424), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n358), .A3(new_n648), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n303), .A2(new_n680), .A3(new_n612), .A4(new_n646), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT97), .B(G146), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G48));
  AND2_X1   g497(.A1(new_n303), .A2(new_n354), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n283), .B1(new_n411), .B2(new_n414), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n423), .A2(KEYINPUT98), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(G469), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n425), .A2(new_n689), .A3(new_n357), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n690), .A2(new_n611), .A3(new_n472), .A4(new_n584), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  AND3_X1   g508(.A1(new_n425), .A2(new_n689), .A3(new_n357), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n303), .A2(new_n354), .A3(new_n695), .A4(new_n624), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  AND4_X1   g511(.A1(new_n357), .A2(new_n425), .A3(new_n689), .A4(new_n589), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n303), .A3(new_n646), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  OAI21_X1  g514(.A(G472), .B1(new_n299), .B2(G902), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n284), .B(KEYINPUT99), .Z(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n279), .A2(new_n265), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n294), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n291), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n701), .A2(new_n354), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n622), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT100), .B1(new_n599), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n711), .B(new_n622), .C1(new_n540), .C2(new_n545), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n690), .A2(new_n472), .A3(new_n584), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n482), .ZN(G24));
  NOR2_X1   g531(.A1(new_n690), .A2(new_n472), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n610), .B(new_n649), .C1(new_n540), .C2(new_n545), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n595), .A2(new_n719), .A3(new_n639), .A4(new_n706), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  NOR2_X1   g536(.A1(new_n415), .A2(new_n416), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT81), .B1(new_n423), .B2(new_n359), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n432), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n357), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT101), .B1(new_n679), .B2(new_n358), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n671), .A2(new_n434), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n719), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n684), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  OR3_X1    g549(.A1(new_n296), .A2(KEYINPUT103), .A3(KEYINPUT32), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT103), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n297), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n354), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n733), .A2(new_n735), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n219), .ZN(G33));
  NAND3_X1  g559(.A1(new_n731), .A2(new_n684), .A3(new_n651), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n430), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n428), .A2(KEYINPUT45), .A3(new_n429), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(G469), .A2(G902), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT104), .A3(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n425), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n357), .A3(new_n655), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n599), .A2(new_n610), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n599), .A2(new_n765), .A3(new_n610), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n596), .A3(new_n639), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT44), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n729), .B(KEYINPUT106), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NOR4_X1   g586(.A1(new_n303), .A2(new_n354), .A3(new_n719), .A4(new_n729), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n357), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT47), .B1(new_n760), .B2(new_n357), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND3_X1  g591(.A1(new_n354), .A2(new_n434), .A3(new_n357), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n425), .A2(new_n689), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n763), .B(new_n778), .C1(new_n779), .C2(KEYINPUT49), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT107), .Z(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT108), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n670), .A3(new_n674), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT109), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n684), .A2(new_n691), .B1(new_n715), .B2(new_n714), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n720), .A2(new_n727), .A3(new_n730), .A4(new_n728), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n622), .A2(new_n648), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n621), .A2(new_n644), .A3(new_n620), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n303), .A2(new_n433), .A3(new_n730), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n696), .A2(new_n699), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n791), .A3(new_n792), .A4(new_n746), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n744), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n472), .B1(new_n710), .B2(new_n712), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n669), .A2(new_n680), .A3(new_n795), .A4(new_n639), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n681), .A3(new_n652), .A4(new_n721), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n473), .A2(new_n480), .A3(new_n585), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n613), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT110), .B1(new_n591), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  OAI221_X1 g617(.A(new_n803), .B1(new_n613), .B2(new_n800), .C1(new_n355), .C2(new_n590), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n600), .A2(new_n709), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n433), .A2(new_n596), .A3(new_n354), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n800), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n640), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n802), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n652), .A2(new_n721), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n794), .A2(new_n799), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n794), .A2(new_n799), .A3(KEYINPUT53), .A4(new_n809), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n802), .A2(new_n804), .A3(new_n808), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n793), .A3(new_n744), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT53), .A4(new_n799), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n774), .B2(new_n775), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n760), .A2(new_n357), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n357), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n425), .A2(new_n689), .A3(new_n358), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n764), .A2(new_n581), .A3(new_n766), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n708), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n770), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n835), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n690), .A2(new_n729), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n701), .A2(new_n644), .A3(new_n707), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n434), .B1(new_n672), .B2(new_n673), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n836), .A3(new_n695), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n836), .A3(KEYINPUT50), .A4(new_n695), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n354), .A2(new_n581), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n600), .A2(new_n610), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n670), .A2(new_n842), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT51), .B1(new_n840), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n843), .A2(new_n739), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT48), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n836), .A2(new_n718), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n670), .A2(new_n842), .A3(new_n612), .A4(new_n852), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(new_n578), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n774), .A2(new_n775), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n838), .B1(new_n868), .B2(new_n833), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n851), .A2(new_n855), .A3(KEYINPUT51), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n861), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n825), .B1(new_n858), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n861), .A2(new_n864), .A3(new_n866), .ZN(new_n873));
  INV_X1    g687(.A(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n833), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n839), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n856), .B1(new_n834), .B2(new_n839), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n877), .B(KEYINPUT118), .C1(KEYINPUT51), .C2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n818), .A2(new_n813), .A3(new_n799), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n821), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n824), .A2(new_n880), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n887), .A2(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n885), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT112), .B1(new_n821), .B2(KEYINPUT54), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT119), .B1(new_n892), .B2(new_n880), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n785), .B1(new_n889), .B2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n883), .A2(new_n283), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n447), .A2(new_n449), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(new_n455), .Z(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n337), .A2(G952), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT121), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n901), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n903), .A2(new_n909), .ZN(G51));
  XNOR2_X1  g724(.A(new_n883), .B(new_n884), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n752), .B(KEYINPUT122), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n411), .B2(new_n414), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n883), .A2(new_n283), .A3(new_n751), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n904), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  INV_X1    g732(.A(new_n618), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n904), .ZN(G60));
  OR2_X1    g736(.A1(new_n606), .A2(new_n607), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n892), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n924), .A2(new_n926), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n906), .B1(new_n911), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(G63));
  INV_X1    g744(.A(new_n883), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n340), .B2(new_n341), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n931), .A2(new_n636), .A3(new_n637), .A4(new_n933), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n905), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n583), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  AND3_X1   g756(.A1(new_n809), .A2(new_n786), .A3(new_n792), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n899), .B1(G898), .B2(new_n337), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G69));
  AND2_X1   g760(.A1(new_n810), .A2(new_n681), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n677), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  INV_X1    g763(.A(new_n776), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n611), .B1(new_n600), .B2(new_n709), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n658), .A2(new_n684), .A3(new_n730), .A4(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n771), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n771), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n270), .ZN(new_n958));
  MUX2_X1   g772(.A(new_n257), .B(new_n958), .S(KEYINPUT30), .Z(new_n959));
  NOR2_X1   g773(.A1(new_n505), .A2(new_n506), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n337), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(G900), .B1(new_n961), .B2(G227), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(G953), .ZN(new_n965));
  INV_X1    g779(.A(new_n746), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n744), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT126), .Z(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n337), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n739), .A2(new_n472), .A3(new_n713), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n762), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT125), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n771), .A2(new_n776), .A3(new_n947), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n969), .A2(new_n974), .B1(G227), .B2(G953), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n963), .B(new_n965), .C1(new_n975), .C2(new_n962), .ZN(G72));
  OAI211_X1 g790(.A(new_n951), .B(new_n943), .C1(new_n956), .C2(new_n955), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT63), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT127), .Z(new_n980));
  AOI22_X1  g794(.A1(new_n977), .A2(new_n980), .B1(new_n258), .B2(new_n259), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n974), .A2(new_n943), .A3(new_n968), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n265), .B1(new_n982), .B2(new_n980), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n267), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n267), .B2(new_n663), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n904), .B1(new_n821), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G57));
endmodule


