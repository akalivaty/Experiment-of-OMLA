

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U325 ( .A(n411), .B(n410), .Z(n293) );
  AND2_X1 U326 ( .A1(n572), .A2(n561), .ZN(n386) );
  INV_X1 U327 ( .A(KEYINPUT122), .ZN(n409) );
  XNOR2_X1 U328 ( .A(n409), .B(KEYINPUT54), .ZN(n410) );
  XNOR2_X1 U329 ( .A(n353), .B(KEYINPUT32), .ZN(n354) );
  XNOR2_X1 U330 ( .A(n355), .B(n354), .ZN(n358) );
  XNOR2_X1 U331 ( .A(n403), .B(n359), .ZN(n360) );
  XNOR2_X1 U332 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U333 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U335 ( .A(KEYINPUT41), .B(n575), .Z(n561) );
  XOR2_X1 U336 ( .A(n330), .B(n329), .Z(n526) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n452) );
  XNOR2_X1 U338 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n295) );
  NAND2_X1 U340 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(KEYINPUT76), .Z(n302) );
  XOR2_X1 U343 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U344 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n336) );
  XOR2_X1 U346 ( .A(KEYINPUT73), .B(G85GAT), .Z(n300) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n356) );
  XNOR2_X1 U349 ( .A(n336), .B(n356), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U351 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n304) );
  XNOR2_X1 U352 ( .A(G134GAT), .B(KEYINPUT64), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U354 ( .A(n306), .B(n305), .Z(n311) );
  XNOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n307), .B(G162GAT), .ZN(n436) );
  XOR2_X1 U357 ( .A(G92GAT), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n399) );
  XNOR2_X1 U360 ( .A(n436), .B(n399), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n554) );
  XNOR2_X1 U362 ( .A(n554), .B(KEYINPUT77), .ZN(n536) );
  XOR2_X1 U363 ( .A(KEYINPUT85), .B(G176GAT), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT84), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n330) );
  XOR2_X1 U366 ( .A(KEYINPUT82), .B(G134GAT), .Z(n315) );
  XNOR2_X1 U367 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(G113GAT), .B(n316), .Z(n425) );
  XOR2_X1 U370 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n318) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n397) );
  XOR2_X1 U373 ( .A(KEYINPUT86), .B(n397), .Z(n320) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n425), .B(n321), .ZN(n328) );
  XOR2_X1 U377 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n323) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G71GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(n324), .B(G190GAT), .Z(n326) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G127GAT), .Z(n375) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(n375), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  INV_X1 U385 ( .A(n526), .ZN(n451) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G113GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(G50GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(n333), .B(G22GAT), .Z(n335) );
  XOR2_X1 U390 ( .A(G1GAT), .B(KEYINPUT69), .Z(n376) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(n376), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U393 ( .A(n336), .B(KEYINPUT29), .Z(n338) );
  NAND2_X1 U394 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(n340), .B(n339), .Z(n348) );
  XOR2_X1 U397 ( .A(KEYINPUT65), .B(KEYINPUT68), .Z(n342) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G197GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U400 ( .A(G8GAT), .B(KEYINPUT67), .Z(n344) );
  XNOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n572) );
  XOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n350) );
  XNOR2_X1 U406 ( .A(G78GAT), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n363) );
  XOR2_X1 U408 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n352) );
  XNOR2_X1 U409 ( .A(G71GAT), .B(G57GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n370) );
  XOR2_X1 U411 ( .A(KEYINPUT72), .B(G148GAT), .Z(n432) );
  XNOR2_X1 U412 ( .A(n370), .B(n432), .ZN(n355) );
  AND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n356), .B(KEYINPUT71), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n361) );
  XOR2_X1 U416 ( .A(G176GAT), .B(G64GAT), .Z(n403) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(G92GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n575) );
  XOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n365) );
  XNOR2_X1 U420 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n380) );
  XOR2_X1 U422 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n367) );
  NAND2_X1 U423 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n368), .B(KEYINPUT79), .Z(n372) );
  XNOR2_X1 U426 ( .A(G22GAT), .B(G155GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n369), .B(G78GAT), .ZN(n442) );
  XNOR2_X1 U428 ( .A(n442), .B(n370), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n374) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(G183GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n373), .B(G211GAT), .ZN(n398) );
  XOR2_X1 U432 ( .A(n374), .B(n398), .Z(n378) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(n380), .B(n379), .Z(n550) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n381) );
  XOR2_X1 U437 ( .A(n536), .B(n381), .Z(n582) );
  NOR2_X1 U438 ( .A1(n550), .A2(n582), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT45), .B(n382), .Z(n383) );
  NOR2_X1 U440 ( .A1(n575), .A2(n383), .ZN(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT114), .B(n384), .Z(n385) );
  NOR2_X1 U442 ( .A1(n572), .A2(n385), .ZN(n393) );
  XNOR2_X1 U443 ( .A(n386), .B(KEYINPUT46), .ZN(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT112), .B(n550), .Z(n564) );
  INV_X1 U445 ( .A(n554), .ZN(n387) );
  OR2_X1 U446 ( .A1(n564), .A2(n387), .ZN(n388) );
  OR2_X1 U447 ( .A1(n389), .A2(n388), .ZN(n391) );
  XOR2_X1 U448 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U450 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(KEYINPUT48), .ZN(n525) );
  XOR2_X1 U452 ( .A(G204GAT), .B(KEYINPUT87), .Z(n396) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n433) );
  XNOR2_X1 U455 ( .A(n397), .B(n433), .ZN(n407) );
  XOR2_X1 U456 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n401) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U459 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n517) );
  XNOR2_X1 U463 ( .A(n517), .B(KEYINPUT121), .ZN(n408) );
  NOR2_X1 U464 ( .A1(n525), .A2(n408), .ZN(n411) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G127GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U471 ( .A(KEYINPUT1), .B(G148GAT), .Z(n417) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G155GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n419), .B(n418), .Z(n427) );
  XOR2_X1 U475 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n421) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n441) );
  XOR2_X1 U478 ( .A(G57GAT), .B(n441), .Z(n423) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n514) );
  INV_X1 U484 ( .A(n514), .ZN(n569) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n431) );
  XNOR2_X1 U486 ( .A(G211GAT), .B(KEYINPUT22), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n446) );
  XOR2_X1 U488 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U489 ( .A(G218GAT), .B(G106GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(n436), .Z(n438) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n464) );
  AND2_X1 U498 ( .A1(n569), .A2(n464), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n293), .A2(n447), .ZN(n449) );
  NOR2_X1 U500 ( .A1(n451), .A2(n450), .ZN(n565) );
  NAND2_X1 U501 ( .A1(n536), .A2(n565), .ZN(n453) );
  INV_X1 U502 ( .A(n572), .ZN(n500) );
  OR2_X1 U503 ( .A1(n500), .A2(n575), .ZN(n486) );
  NAND2_X1 U504 ( .A1(n526), .A2(n517), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n464), .A2(n454), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT25), .ZN(n459) );
  NOR2_X1 U507 ( .A1(n526), .A2(n464), .ZN(n457) );
  XNOR2_X1 U508 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n456) );
  XOR2_X1 U509 ( .A(n457), .B(n456), .Z(n571) );
  XNOR2_X1 U510 ( .A(n517), .B(KEYINPUT27), .ZN(n462) );
  AND2_X1 U511 ( .A1(n571), .A2(n462), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT96), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n514), .A2(n461), .ZN(n468) );
  NAND2_X1 U515 ( .A1(n462), .A2(n514), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT93), .ZN(n541) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n464), .Z(n520) );
  INV_X1 U518 ( .A(n520), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n541), .A2(n465), .ZN(n528) );
  NOR2_X1 U520 ( .A1(n526), .A2(n528), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT94), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n483) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n470) );
  OR2_X1 U524 ( .A1(n536), .A2(n550), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(n471) );
  OR2_X1 U526 ( .A1(n483), .A2(n471), .ZN(n501) );
  NOR2_X1 U527 ( .A1(n486), .A2(n501), .ZN(n480) );
  NAND2_X1 U528 ( .A1(n480), .A2(n514), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT34), .B(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT97), .Z(n475) );
  NAND2_X1 U532 ( .A1(n480), .A2(n517), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U535 ( .A1(n480), .A2(n526), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT98), .Z(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n520), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT100), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NOR2_X1 U543 ( .A1(n483), .A2(n582), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n550), .A2(n484), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n485), .Z(n513) );
  NOR2_X1 U546 ( .A1(n513), .A2(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n495), .A2(n514), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  XOR2_X1 U551 ( .A(G36GAT), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U552 ( .A1(n495), .A2(n517), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n526), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n520), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n499) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n500), .A2(n561), .ZN(n512) );
  OR2_X1 U564 ( .A1(n501), .A2(n512), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT106), .B(n502), .Z(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n514), .ZN(n503) );
  XOR2_X1 U567 ( .A(n504), .B(n503), .Z(G1332GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n517), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n507), .A2(n526), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U573 ( .A1(n507), .A2(n520), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT108), .Z(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT110), .B(n515), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n526), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT115), .Z(n530) );
  INV_X1 U590 ( .A(n525), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n526), .A2(n542), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n572), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n532) );
  NAND2_X1 U596 ( .A1(n537), .A2(n561), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n564), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  AND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n571), .A2(n543), .ZN(n553) );
  INV_X1 U608 ( .A(n553), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n551), .A2(n572), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(n547), .Z(n549) );
  NAND2_X1 U615 ( .A1(n551), .A2(n561), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  INV_X1 U617 ( .A(n550), .ZN(n579) );
  NAND2_X1 U618 ( .A1(n579), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT120), .B(n555), .Z(n556) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n565), .A2(n572), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT59), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(n568), .Z(n574) );
  AND2_X1 U636 ( .A1(n293), .A2(n569), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n581) );
  INV_X1 U638 ( .A(n581), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n578), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

