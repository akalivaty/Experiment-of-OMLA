//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G952), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n189), .B1(G234), .B2(G237), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT21), .B(G898), .Z(new_n192));
  NAND2_X1  g006(.A1(G234), .A2(G237), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n193), .A2(G902), .A3(G953), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n192), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G210), .B1(G237), .B2(G902), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(G104), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT81), .A3(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(G116), .A2(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G119), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G113), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n216), .A2(new_n217), .B1(new_n211), .B2(new_n212), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(KEYINPUT3), .C1(new_n202), .C2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n202), .A2(G107), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT79), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n201), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(KEYINPUT79), .B2(new_n227), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(KEYINPUT79), .A2(new_n227), .B1(new_n199), .B2(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n227), .A2(KEYINPUT79), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n223), .B(new_n224), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT80), .B1(new_n236), .B2(G101), .ZN(new_n237));
  AOI211_X1 g051(.A(new_n206), .B(new_n221), .C1(new_n233), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n239), .A3(G101), .ZN(new_n240));
  INV_X1    g054(.A(new_n213), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n207), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n214), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(new_n233), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n239), .B1(new_n236), .B2(G101), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G110), .B(G122), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n238), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n257), .A3(new_n259), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n256), .A2(KEYINPUT1), .A3(G146), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(new_n268), .C1(G128), .C2(new_n253), .ZN(new_n269));
  INV_X1    g083(.A(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n188), .A2(G224), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT86), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n271), .A4(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n213), .A2(KEYINPUT5), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n214), .B1(new_n279), .B2(new_n219), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n235), .B1(new_n201), .B2(new_n228), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n225), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n231), .B1(new_n282), .B2(new_n232), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n236), .A2(KEYINPUT80), .A3(G101), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n205), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT8), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n250), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n221), .B1(new_n245), .B2(new_n205), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n251), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n278), .B(KEYINPUT87), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n250), .B1(new_n238), .B2(new_n247), .ZN(new_n295));
  INV_X1    g109(.A(new_n221), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n245), .A2(new_n205), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n250), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT4), .B1(new_n282), .B2(new_n232), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n233), .B2(new_n237), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n298), .C1(new_n300), .C2(new_n244), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(KEYINPUT6), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(new_n250), .C1(new_n238), .C2(new_n247), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n272), .B(new_n274), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n197), .B1(new_n294), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n290), .A2(new_n291), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n301), .A3(new_n293), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n308), .A2(new_n310), .A3(new_n306), .A4(new_n197), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n187), .B(new_n196), .C1(new_n307), .C2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n313), .A2(new_n314), .A3(G953), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n256), .A2(G128), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n256), .B2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n265), .A2(KEYINPUT92), .A3(G143), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n318), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n324));
  INV_X1    g138(.A(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G122), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G116), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n209), .A2(G122), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  XNOR2_X1  g146(.A(G116), .B(G122), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n199), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n321), .A2(new_n322), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n317), .A3(new_n319), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT14), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n329), .A2(new_n330), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G107), .B1(new_n330), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n334), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n319), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G134), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n337), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n316), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n323), .A2(new_n326), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G134), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n325), .B1(new_n321), .B2(new_n322), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n350), .A2(new_n317), .B1(new_n332), .B2(new_n334), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n337), .ZN(new_n353));
  INV_X1    g167(.A(new_n343), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n355), .A3(new_n315), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n347), .A2(new_n356), .A3(KEYINPUT93), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT93), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n359), .B(new_n316), .C1(new_n339), .C2(new_n346), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n308), .A4(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G478), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT15), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n361), .A2(new_n363), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT89), .ZN(new_n369));
  XNOR2_X1  g183(.A(G113), .B(G122), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(new_n202), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G125), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(KEYINPUT74), .A3(G125), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  OAI211_X1 g195(.A(G146), .B(new_n375), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(G237), .A2(G953), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G143), .A3(G214), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(G143), .B1(new_n383), .B2(G214), .ZN(new_n386));
  OAI21_X1  g200(.A(G131), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(G131), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n270), .A2(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n373), .A2(new_n395), .A3(new_n378), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n376), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT19), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n379), .A2(new_n398), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n393), .A2(new_n399), .A3(new_n258), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n388), .A2(new_n384), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT18), .A3(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n258), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n397), .B2(new_n258), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n388), .A2(new_n384), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n371), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n387), .A2(new_n390), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n381), .B1(new_n396), .B2(new_n376), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n258), .B1(new_n413), .B2(new_n374), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n403), .A2(KEYINPUT17), .A3(G131), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n382), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n416), .A2(new_n371), .A3(new_n409), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n369), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n371), .A3(new_n409), .ZN(new_n420));
  INV_X1    g234(.A(new_n409), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n392), .B2(new_n401), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n371), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n369), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n371), .B1(new_n416), .B2(new_n409), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n308), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT90), .B(G475), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n419), .A2(new_n425), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n367), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n312), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n383), .A2(G210), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT27), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT26), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n435), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT26), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n437), .A2(new_n441), .A3(G101), .ZN(new_n442));
  AOI21_X1  g256(.A(G101), .B1(new_n437), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n445));
  INV_X1    g259(.A(new_n243), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n268), .B1(new_n253), .B2(G128), .ZN(new_n447));
  INV_X1    g261(.A(new_n267), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT11), .B1(new_n317), .B2(G137), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT65), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n452), .B2(G134), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n317), .A2(KEYINPUT65), .A3(G137), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(new_n458), .A3(new_n389), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n452), .A2(G134), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n317), .A2(G137), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n389), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n449), .B1(new_n464), .B2(KEYINPUT67), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n450), .A2(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n462), .B1(new_n466), .B2(new_n389), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n458), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT66), .A2(G131), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n454), .A2(new_n458), .A3(KEYINPUT66), .A4(G131), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n263), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n446), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n269), .A2(new_n463), .A3(new_n459), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(new_n446), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n445), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n446), .A3(new_n477), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n444), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n473), .A2(new_n474), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n465), .A2(new_n469), .B1(new_n485), .B2(new_n263), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n243), .B(new_n484), .C1(new_n486), .C2(KEYINPUT30), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n478), .A2(new_n442), .A3(new_n443), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n489), .A3(new_n488), .A4(KEYINPUT31), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n434), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n483), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n444), .A2(new_n480), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n269), .B1(new_n467), .B2(new_n468), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n475), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n499), .B1(new_n505), .B2(new_n243), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT31), .B1(new_n506), .B2(new_n488), .ZN(new_n507));
  INV_X1    g321(.A(new_n493), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n498), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT32), .A3(new_n495), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n487), .A2(new_n480), .ZN(new_n511));
  INV_X1    g325(.A(new_n444), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT29), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n479), .A2(new_n444), .A3(new_n482), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n480), .A2(KEYINPUT71), .A3(new_n481), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT71), .B1(new_n480), .B2(new_n481), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n444), .A2(KEYINPUT29), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n475), .A2(new_n477), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n243), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n480), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT70), .B1(new_n522), .B2(KEYINPUT28), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n446), .B1(new_n475), .B2(new_n477), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n478), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n518), .B(new_n519), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT28), .B1(new_n478), .B2(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n525), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n518), .A4(new_n519), .ZN(new_n534));
  AOI221_X4 g348(.A(G902), .B1(new_n513), .B2(new_n514), .C1(new_n528), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G472), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n497), .B(new_n510), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G469), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT83), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n188), .A2(G227), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(G140), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT78), .B(G110), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n205), .B1(new_n447), .B2(new_n448), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n283), .B2(new_n284), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT82), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n547), .B1(new_n237), .B2(new_n233), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(KEYINPUT10), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n485), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n245), .A2(new_n246), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n240), .A2(new_n263), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n557), .A2(new_n558), .B1(new_n553), .B2(KEYINPUT10), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n556), .B1(new_n555), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n546), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT82), .B1(new_n549), .B2(new_n550), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n553), .A2(new_n552), .A3(KEYINPUT10), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n559), .B(new_n556), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n269), .B1(new_n245), .B2(new_n205), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n485), .B1(new_n566), .B2(new_n553), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT12), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n569), .B(new_n485), .C1(new_n566), .C2(new_n553), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n545), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n541), .B1(new_n562), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n559), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n485), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n565), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT83), .B1(new_n575), .B2(new_n546), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n540), .B(new_n308), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n546), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n565), .A3(new_n545), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(G469), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n540), .A2(new_n308), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n539), .B1(new_n577), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n265), .A2(G119), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n210), .A2(G128), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT24), .B(G110), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n210), .B2(G128), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT23), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT23), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n595), .A3(new_n587), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n590), .B1(new_n596), .B2(G110), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n382), .A2(new_n597), .A3(new_n405), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT75), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n382), .A2(new_n597), .A3(new_n600), .A4(new_n405), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n382), .A2(new_n414), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n588), .A2(new_n589), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n596), .B2(G110), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT22), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n452), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n612), .A3(G137), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(new_n599), .A3(new_n601), .A4(new_n605), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n314), .B1(G234), .B2(new_n308), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(new_n622), .B2(G902), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n619), .A2(new_n621), .A3(KEYINPUT25), .A4(new_n308), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(KEYINPUT77), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n624), .B1(new_n628), .B2(KEYINPUT77), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n433), .A2(new_n537), .A3(new_n585), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  OAI21_X1  g449(.A(G472), .B1(new_n494), .B2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n509), .A2(new_n495), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n585), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT95), .Z(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n357), .A2(new_n642), .A3(new_n360), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n347), .A2(new_n356), .A3(KEYINPUT33), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n362), .A2(G902), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n357), .A2(new_n308), .A3(new_n360), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n362), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(KEYINPUT96), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT96), .B1(new_n646), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n312), .A2(new_n431), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n641), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n417), .A2(new_n426), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n430), .B1(new_n659), .B2(G902), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n419), .A2(new_n425), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(KEYINPUT97), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n365), .A2(new_n366), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n419), .A2(new_n665), .A3(new_n425), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n658), .B1(new_n312), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n418), .A2(KEYINPUT20), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n424), .B1(new_n423), .B2(new_n369), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT97), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n660), .A3(new_n666), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n367), .ZN(new_n673));
  INV_X1    g487(.A(new_n187), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n310), .A2(new_n306), .A3(new_n308), .ZN(new_n675));
  INV_X1    g489(.A(new_n197), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n294), .A2(new_n197), .A3(new_n306), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n679), .A3(KEYINPUT98), .A4(new_n196), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n641), .B1(new_n668), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NOR2_X1   g497(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n606), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n625), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n630), .B2(new_n631), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n433), .A2(new_n585), .A3(new_n639), .A4(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  OAI21_X1  g504(.A(new_n187), .B1(new_n307), .B2(new_n311), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n195), .B2(G900), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n194), .A2(KEYINPUT99), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n191), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n663), .A2(new_n664), .A3(new_n666), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n537), .A2(new_n585), .A3(new_n698), .A4(new_n687), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n687), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT32), .B1(new_n509), .B2(new_n495), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n494), .A2(new_n434), .A3(new_n496), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n528), .A2(new_n534), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n513), .A2(new_n514), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n308), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G472), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n702), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(KEYINPUT100), .A3(new_n585), .A4(new_n698), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XOR2_X1   g527(.A(new_n696), .B(KEYINPUT103), .Z(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(KEYINPUT39), .Z(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n585), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n677), .A2(new_n678), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT38), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n187), .B1(new_n365), .B2(new_n366), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n431), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n720), .A2(new_n702), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n512), .B1(new_n487), .B2(new_n480), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n308), .B1(new_n522), .B2(new_n444), .ZN(new_n725));
  OAI21_X1  g539(.A(G472), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n705), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT101), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n705), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n723), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n723), .B2(new_n731), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n718), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  OAI21_X1  g550(.A(new_n660), .B1(new_n669), .B2(new_n670), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n696), .C1(new_n650), .C2(new_n651), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT104), .B1(new_n739), .B2(new_n679), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n691), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n710), .B(new_n585), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  OAI21_X1  g558(.A(new_n308), .B1(new_n572), .B2(new_n576), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G469), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n746), .A2(new_n538), .A3(new_n577), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n632), .B1(new_n705), .B2(new_n709), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n653), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND2_X1  g565(.A1(new_n668), .A2(new_n680), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n748), .A3(new_n747), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  NAND4_X1  g568(.A1(new_n747), .A2(new_n537), .A3(new_n433), .A4(new_n687), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n719), .A2(new_n722), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT105), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n719), .A2(new_n722), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n517), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n515), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n531), .B2(new_n525), .ZN(new_n764));
  OAI22_X1  g578(.A1(new_n507), .A2(new_n508), .B1(new_n764), .B2(new_n444), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n495), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n633), .A2(new_n636), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n747), .A2(new_n761), .A3(new_n767), .A4(new_n196), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND3_X1  g583(.A1(new_n687), .A2(new_n636), .A3(new_n766), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n738), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n747), .A2(new_n679), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NAND2_X1  g587(.A1(new_n579), .A2(new_n580), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n580), .A2(KEYINPUT106), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(G469), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n577), .A3(new_n583), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n719), .A2(new_n674), .A3(new_n539), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n748), .A2(new_n739), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n510), .A2(new_n497), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n783), .A2(KEYINPUT107), .B1(G472), .B2(new_n708), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n705), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n632), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n738), .A2(new_n782), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n779), .A2(new_n780), .A3(new_n788), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n781), .A2(new_n782), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n389), .ZN(G33));
  INV_X1    g605(.A(new_n697), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n748), .A2(new_n792), .A3(new_n779), .A4(new_n780), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  AOI21_X1  g608(.A(KEYINPUT106), .B1(new_n579), .B2(new_n580), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n580), .A2(KEYINPUT106), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT45), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n540), .B1(new_n774), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n582), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n577), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(KEYINPUT108), .A3(new_n538), .A4(new_n716), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n538), .B1(new_n802), .B2(new_n803), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n715), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT43), .B1(new_n652), .B2(new_n737), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n646), .A2(new_n648), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n649), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT43), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n431), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n809), .A2(new_n638), .A3(new_n687), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n677), .A2(new_n678), .A3(new_n187), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n805), .A2(new_n808), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G137), .ZN(G39));
  NAND2_X1  g637(.A1(new_n807), .A2(KEYINPUT47), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n538), .C1(new_n802), .C2(new_n803), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n537), .A2(new_n633), .A3(new_n738), .A4(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND2_X1  g643(.A1(new_n746), .A2(new_n577), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT110), .Z(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT49), .ZN(new_n832));
  INV_X1    g646(.A(new_n731), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n633), .A2(new_n187), .A3(new_n538), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT109), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n720), .A2(new_n737), .A3(new_n652), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n633), .A2(new_n636), .A3(new_n766), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n809), .A2(new_n190), .A3(new_n815), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n809), .A2(KEYINPUT114), .A3(new_n190), .A4(new_n815), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n679), .A3(new_n747), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n846), .A3(new_n679), .A4(new_n747), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n820), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n747), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n841), .B2(new_n842), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n787), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n841), .A2(new_n842), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n747), .A3(new_n787), .A4(new_n849), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n852), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n633), .A2(new_n190), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n731), .A2(new_n850), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n652), .A2(new_n431), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n189), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n848), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n824), .A2(new_n826), .B1(new_n539), .B2(new_n831), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n843), .A2(new_n849), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n720), .A2(new_n187), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n843), .A2(new_n747), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT50), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(KEYINPUT50), .ZN(new_n870));
  INV_X1    g684(.A(new_n770), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n851), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n813), .A2(new_n737), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n869), .A2(new_n870), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n863), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n872), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n869), .A4(new_n870), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n864), .A2(new_n865), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n701), .A2(new_n711), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n696), .A2(new_n538), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n686), .B(new_n886), .C1(new_n630), .C2(new_n631), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n582), .B1(new_n797), .B2(G469), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n577), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n761), .A3(new_n727), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n743), .A2(new_n890), .A3(new_n772), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n885), .A2(new_n891), .A3(KEYINPUT52), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n743), .A2(new_n890), .A3(new_n772), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n712), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n367), .A2(new_n696), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n672), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n849), .A2(KEYINPUT112), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT112), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n663), .A2(new_n367), .A3(new_n666), .A4(new_n696), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n820), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n710), .A2(new_n585), .A3(new_n899), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n771), .A2(new_n779), .A3(new_n780), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n793), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n790), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n812), .A2(new_n737), .A3(new_n649), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n432), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n312), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n585), .A3(new_n633), .A4(new_n639), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n634), .A2(new_n688), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT111), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n634), .A2(new_n688), .A3(new_n910), .A4(KEYINPUT111), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND4_X1   g729(.A1(new_n749), .A2(new_n753), .A3(new_n768), .A4(new_n755), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n906), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n896), .A2(new_n917), .A3(KEYINPUT53), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT52), .B1(new_n885), .B2(new_n891), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n894), .A2(new_n893), .A3(new_n712), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n906), .A2(new_n915), .A3(new_n916), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n896), .B2(new_n917), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n922), .A2(new_n923), .A3(new_n919), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n884), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n837), .B1(new_n930), .B2(new_n931), .ZN(G75));
  NAND2_X1  g746(.A1(new_n918), .A2(new_n924), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(G210), .A3(G902), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n302), .A2(new_n304), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n305), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n934), .B2(new_n936), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n188), .A2(G952), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(new_n582), .B(KEYINPUT57), .ZN(new_n944));
  INV_X1    g758(.A(new_n926), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n925), .B1(new_n918), .B2(new_n924), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n572), .A2(new_n576), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n933), .A2(G902), .A3(new_n798), .A4(new_n800), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G54));
  INV_X1    g765(.A(new_n942), .ZN(new_n952));
  NAND2_X1  g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT119), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n308), .B(new_n955), .C1(new_n918), .C2(new_n924), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n423), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n933), .A2(G902), .A3(new_n423), .A4(new_n954), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT120), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT120), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G60));
  XNOR2_X1  g775(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n362), .A2(new_n308), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n929), .B2(new_n926), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n643), .A2(new_n644), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n952), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n966), .B(new_n964), .C1(new_n929), .C2(new_n926), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT122), .Z(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT60), .Z(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n927), .B2(new_n928), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n942), .B1(new_n974), .B2(new_n622), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n918), .B2(new_n924), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n685), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n975), .B(new_n978), .C1(new_n979), .C2(KEYINPUT61), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(new_n952), .C1(new_n977), .C2(new_n623), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n952), .B1(new_n977), .B2(new_n623), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n933), .A2(new_n685), .A3(new_n973), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n981), .B(new_n982), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n985), .ZN(G66));
  NAND3_X1  g800(.A1(new_n192), .A2(G224), .A3(G953), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n915), .A2(new_n916), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n937), .B1(G898), .B2(new_n188), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(G69));
  AND3_X1   g805(.A1(new_n712), .A2(new_n743), .A3(new_n772), .ZN(new_n992));
  INV_X1    g806(.A(new_n793), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n790), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n828), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n787), .A2(new_n761), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n805), .B(new_n808), .C1(new_n821), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n188), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n505), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n694), .B2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT124), .ZN(new_n1003));
  INV_X1    g817(.A(G227), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n1004), .B2(new_n694), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n999), .A2(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n735), .A2(new_n992), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n908), .A2(new_n820), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n717), .A2(new_n748), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1009), .A2(new_n822), .A3(new_n828), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n735), .B2(new_n992), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n188), .B(new_n1001), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1006), .A2(new_n1007), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1007), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1015), .A2(new_n1016), .ZN(G72));
  NOR3_X1   g831(.A1(new_n1012), .A2(new_n988), .A3(new_n1013), .ZN(new_n1018));
  XNOR2_X1  g832(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n536), .A2(new_n308), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n724), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT127), .B1(new_n511), .B2(new_n512), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1023), .A2(new_n506), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n511), .A2(KEYINPUT127), .A3(new_n512), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n933), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n511), .A2(new_n444), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n995), .A2(new_n915), .A3(new_n916), .A4(new_n997), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1021), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(KEYINPUT126), .B1(new_n1033), .B2(new_n942), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT126), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1035), .B(new_n952), .C1(new_n1036), .C2(new_n1030), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1028), .B1(new_n1034), .B2(new_n1037), .ZN(G57));
endmodule


