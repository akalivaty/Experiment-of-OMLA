

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770;

  NAND2_X1 U372 ( .A1(n404), .A2(n402), .ZN(n375) );
  NOR2_X2 U373 ( .A1(n653), .A2(n654), .ZN(n651) );
  INV_X1 U374 ( .A(G953), .ZN(n759) );
  NAND2_X2 U375 ( .A1(n421), .A2(n420), .ZN(n419) );
  XNOR2_X2 U376 ( .A(n533), .B(KEYINPUT0), .ZN(n430) );
  NOR2_X2 U377 ( .A1(n690), .A2(n599), .ZN(n639) );
  XNOR2_X2 U378 ( .A(n395), .B(n394), .ZN(n767) );
  AND2_X2 U379 ( .A1(n604), .A2(n631), .ZN(n395) );
  XNOR2_X2 U380 ( .A(n753), .B(n466), .ZN(n537) );
  AND2_X1 U381 ( .A1(n454), .A2(KEYINPUT2), .ZN(n408) );
  NAND2_X1 U382 ( .A1(n393), .A2(n388), .ZN(n758) );
  XNOR2_X1 U383 ( .A(n389), .B(n363), .ZN(n388) );
  NAND2_X1 U384 ( .A1(n391), .A2(n390), .ZN(n389) );
  XNOR2_X1 U385 ( .A(n444), .B(n362), .ZN(n390) );
  XNOR2_X1 U386 ( .A(n575), .B(KEYINPUT103), .ZN(n607) );
  AND2_X1 U387 ( .A1(n767), .A2(n432), .ZN(n393) );
  INV_X1 U388 ( .A(n712), .ZN(n432) );
  AND2_X1 U389 ( .A1(n441), .A2(n440), .ZN(n411) );
  NAND2_X1 U390 ( .A1(n439), .A2(n359), .ZN(n438) );
  XNOR2_X1 U391 ( .A(n612), .B(n437), .ZN(n598) );
  XNOR2_X1 U392 ( .A(n383), .B(KEYINPUT18), .ZN(n449) );
  XNOR2_X1 U393 ( .A(n494), .B(n369), .ZN(n545) );
  XNOR2_X1 U394 ( .A(n512), .B(n450), .ZN(n535) );
  XNOR2_X1 U395 ( .A(G137), .B(G101), .ZN(n482) );
  INV_X1 U396 ( .A(n573), .ZN(n351) );
  BUF_X1 U397 ( .A(n766), .Z(n352) );
  BUF_X1 U398 ( .A(n624), .Z(n353) );
  NAND2_X2 U399 ( .A1(n422), .A2(n419), .ZN(n376) );
  NAND2_X1 U400 ( .A1(n459), .A2(n586), .ZN(n457) );
  NOR2_X1 U401 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U402 ( .A(G137), .B(G140), .ZN(n540) );
  NOR2_X1 U403 ( .A1(n721), .A2(G902), .ZN(n539) );
  OR2_X1 U404 ( .A1(n737), .A2(G902), .ZN(n474) );
  INV_X1 U405 ( .A(G146), .ZN(n466) );
  INV_X1 U406 ( .A(G110), .ZN(n450) );
  XNOR2_X1 U407 ( .A(n579), .B(KEYINPUT108), .ZN(n427) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(G902), .ZN(n642) );
  XNOR2_X1 U409 ( .A(n463), .B(n392), .ZN(n391) );
  INV_X1 U410 ( .A(KEYINPUT70), .ZN(n392) );
  XOR2_X1 U411 ( .A(G134), .B(G122), .Z(n489) );
  XNOR2_X1 U412 ( .A(G107), .B(G116), .ZN(n488) );
  XOR2_X1 U413 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n491) );
  XNOR2_X1 U414 ( .A(n509), .B(n447), .ZN(n569) );
  XNOR2_X1 U415 ( .A(KEYINPUT13), .B(G475), .ZN(n447) );
  XNOR2_X1 U416 ( .A(n615), .B(KEYINPUT1), .ZN(n564) );
  NAND2_X1 U417 ( .A1(n545), .A2(G221), .ZN(n368) );
  XNOR2_X1 U418 ( .A(n515), .B(n473), .ZN(n754) );
  INV_X1 U419 ( .A(KEYINPUT10), .ZN(n473) );
  NOR2_X1 U420 ( .A1(KEYINPUT2), .A2(n399), .ZN(n398) );
  NAND2_X1 U421 ( .A1(n400), .A2(n472), .ZN(n407) );
  NOR2_X1 U422 ( .A1(n643), .A2(KEYINPUT2), .ZN(n680) );
  INV_X1 U423 ( .A(KEYINPUT78), .ZN(n387) );
  XNOR2_X1 U424 ( .A(n436), .B(n435), .ZN(n599) );
  INV_X1 U425 ( .A(KEYINPUT110), .ZN(n435) );
  NOR2_X1 U426 ( .A1(n598), .A2(n613), .ZN(n436) );
  XNOR2_X1 U427 ( .A(n606), .B(n361), .ZN(n364) );
  AND2_X1 U428 ( .A1(n607), .A2(n605), .ZN(n365) );
  BUF_X1 U429 ( .A(n564), .Z(n650) );
  XNOR2_X1 U430 ( .A(n756), .B(n475), .ZN(n534) );
  XOR2_X1 U431 ( .A(KEYINPUT89), .B(n646), .Z(n736) );
  OR2_X1 U432 ( .A1(G902), .A2(G237), .ZN(n524) );
  XOR2_X1 U433 ( .A(KEYINPUT104), .B(KEYINPUT5), .Z(n480) );
  XNOR2_X1 U434 ( .A(n413), .B(G146), .ZN(n515) );
  INV_X1 U435 ( .A(G125), .ZN(n413) );
  XNOR2_X1 U436 ( .A(n429), .B(n467), .ZN(n753) );
  XNOR2_X1 U437 ( .A(n478), .B(G131), .ZN(n467) );
  XOR2_X1 U438 ( .A(KEYINPUT69), .B(G134), .Z(n478) );
  INV_X1 U439 ( .A(KEYINPUT65), .ZN(n399) );
  INV_X1 U440 ( .A(n642), .ZN(n471) );
  XNOR2_X1 U441 ( .A(n515), .B(n461), .ZN(n518) );
  XNOR2_X1 U442 ( .A(n516), .B(KEYINPUT17), .ZN(n461) );
  INV_X1 U443 ( .A(KEYINPUT91), .ZN(n516) );
  NAND2_X1 U444 ( .A1(G237), .A2(G234), .ZN(n526) );
  INV_X1 U445 ( .A(KEYINPUT86), .ZN(n442) );
  NAND2_X1 U446 ( .A1(n665), .A2(n442), .ZN(n440) );
  NOR2_X1 U447 ( .A1(n654), .A2(n417), .ZN(n416) );
  INV_X1 U448 ( .A(KEYINPUT6), .ZN(n437) );
  XNOR2_X1 U449 ( .A(n543), .B(n371), .ZN(n370) );
  XNOR2_X1 U450 ( .A(n540), .B(KEYINPUT23), .ZN(n371) );
  INV_X1 U451 ( .A(KEYINPUT8), .ZN(n369) );
  XNOR2_X1 U452 ( .A(KEYINPUT7), .B(KEYINPUT105), .ZN(n490) );
  INV_X1 U453 ( .A(KEYINPUT39), .ZN(n443) );
  NOR2_X1 U454 ( .A1(n629), .A2(n664), .ZN(n609) );
  NAND2_X1 U455 ( .A1(n415), .A2(n414), .ZN(n626) );
  INV_X1 U456 ( .A(n623), .ZN(n415) );
  NAND2_X1 U457 ( .A1(n374), .A2(n372), .ZN(n459) );
  NOR2_X1 U458 ( .A1(n650), .A2(n373), .ZN(n372) );
  XNOR2_X1 U459 ( .A(n514), .B(n535), .ZN(n743) );
  XNOR2_X1 U460 ( .A(n544), .B(n367), .ZN(n737) );
  XNOR2_X1 U461 ( .A(n754), .B(n418), .ZN(n544) );
  XNOR2_X1 U462 ( .A(n370), .B(n368), .ZN(n367) );
  XNOR2_X1 U463 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n727), .B(KEYINPUT59), .ZN(n728) );
  XNOR2_X1 U465 ( .A(n682), .B(KEYINPUT80), .ZN(n453) );
  XNOR2_X1 U466 ( .A(n680), .B(n387), .ZN(n386) );
  NOR2_X1 U467 ( .A1(n684), .A2(G953), .ZN(n452) );
  INV_X1 U468 ( .A(KEYINPUT112), .ZN(n394) );
  NAND2_X1 U469 ( .A1(n433), .A2(n650), .ZN(n465) );
  XNOR2_X1 U470 ( .A(n434), .B(KEYINPUT36), .ZN(n433) );
  NAND2_X1 U471 ( .A1(n358), .A2(n365), .ZN(n700) );
  INV_X1 U472 ( .A(n459), .ZN(n696) );
  AND2_X1 U473 ( .A1(n568), .A2(n409), .ZN(n689) );
  NOR2_X1 U474 ( .A1(n650), .A2(n410), .ZN(n409) );
  INV_X1 U475 ( .A(n581), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U477 ( .A(n721), .B(n722), .ZN(n723) );
  AND2_X1 U478 ( .A1(n580), .A2(n456), .ZN(n354) );
  XNOR2_X1 U479 ( .A(G122), .B(KEYINPUT16), .ZN(n355) );
  XOR2_X1 U480 ( .A(G140), .B(G143), .Z(n356) );
  NOR2_X1 U481 ( .A1(n768), .A2(n696), .ZN(n357) );
  AND2_X1 U482 ( .A1(n364), .A2(n632), .ZN(n358) );
  NOR2_X1 U483 ( .A1(n665), .A2(n442), .ZN(n359) );
  INV_X1 U484 ( .A(n605), .ZN(n417) );
  AND2_X1 U485 ( .A1(n685), .A2(n452), .ZN(n360) );
  INV_X1 U486 ( .A(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U487 ( .A(KEYINPUT113), .B(KEYINPUT30), .ZN(n361) );
  INV_X1 U488 ( .A(n626), .ZN(n468) );
  XNOR2_X1 U489 ( .A(n537), .B(n536), .ZN(n721) );
  XNOR2_X1 U490 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n362) );
  XNOR2_X1 U491 ( .A(n641), .B(KEYINPUT82), .ZN(n363) );
  NAND2_X1 U492 ( .A1(n365), .A2(n364), .ZN(n629) );
  NAND2_X1 U493 ( .A1(n366), .A2(KEYINPUT45), .ZN(n425) );
  NAND2_X1 U494 ( .A1(n428), .A2(n427), .ZN(n366) );
  INV_X1 U495 ( .A(n366), .ZN(n421) );
  NOR2_X1 U496 ( .A1(n612), .A2(n613), .ZN(n614) );
  NAND2_X1 U497 ( .A1(n416), .A2(n653), .ZN(n613) );
  NAND2_X1 U498 ( .A1(n612), .A2(n653), .ZN(n373) );
  INV_X1 U499 ( .A(n585), .ZN(n374) );
  XNOR2_X2 U500 ( .A(n451), .B(KEYINPUT22), .ZN(n585) );
  AND2_X1 U501 ( .A1(n426), .A2(n354), .ZN(n420) );
  BUF_X1 U502 ( .A(n498), .Z(n377) );
  NAND2_X1 U503 ( .A1(n422), .A2(n419), .ZN(n455) );
  NAND2_X2 U504 ( .A1(n403), .A2(n407), .ZN(n402) );
  NAND2_X1 U505 ( .A1(n376), .A2(n408), .ZN(n378) );
  NAND2_X1 U506 ( .A1(n455), .A2(n408), .ZN(n681) );
  NAND2_X1 U507 ( .A1(n404), .A2(n402), .ZN(n379) );
  NAND2_X1 U508 ( .A1(n404), .A2(n402), .ZN(n462) );
  XOR2_X1 U509 ( .A(n553), .B(KEYINPUT62), .Z(n645) );
  INV_X1 U510 ( .A(n469), .ZN(n396) );
  NAND2_X1 U511 ( .A1(n498), .A2(n477), .ZN(n381) );
  NAND2_X1 U512 ( .A1(n380), .A2(KEYINPUT4), .ZN(n382) );
  NAND2_X1 U513 ( .A1(n381), .A2(n382), .ZN(n383) );
  INV_X1 U514 ( .A(n498), .ZN(n380) );
  XNOR2_X1 U515 ( .A(n498), .B(n477), .ZN(n429) );
  INV_X1 U516 ( .A(n353), .ZN(n414) );
  XNOR2_X1 U517 ( .A(n448), .B(n743), .ZN(n715) );
  XNOR2_X1 U518 ( .A(n449), .B(n519), .ZN(n448) );
  NAND2_X1 U519 ( .A1(n386), .A2(n378), .ZN(n682) );
  NAND2_X1 U520 ( .A1(n400), .A2(n398), .ZN(n406) );
  AND2_X1 U521 ( .A1(n455), .A2(n454), .ZN(n643) );
  BUF_X1 U522 ( .A(n715), .Z(n384) );
  XNOR2_X1 U523 ( .A(n431), .B(KEYINPUT19), .ZN(n624) );
  BUF_X1 U524 ( .A(n603), .Z(n631) );
  NAND2_X1 U525 ( .A1(n385), .A2(n740), .ZN(n649) );
  XNOR2_X1 U526 ( .A(n644), .B(n645), .ZN(n385) );
  AND2_X2 U527 ( .A1(n405), .A2(n406), .ZN(n404) );
  NAND2_X1 U528 ( .A1(n453), .A2(n360), .ZN(n688) );
  NAND2_X1 U529 ( .A1(n681), .A2(n396), .ZN(n401) );
  AND2_X1 U530 ( .A1(n378), .A2(n397), .ZN(n403) );
  NOR2_X1 U531 ( .A1(n469), .A2(KEYINPUT65), .ZN(n397) );
  INV_X1 U532 ( .A(n376), .ZN(n400) );
  NAND2_X1 U533 ( .A1(n401), .A2(KEYINPUT65), .ZN(n405) );
  AND2_X2 U534 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X2 U535 ( .A(n584), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U536 ( .A1(n411), .A2(n438), .ZN(n431) );
  NAND2_X1 U537 ( .A1(n412), .A2(n557), .ZN(n559) );
  XNOR2_X1 U538 ( .A(n556), .B(KEYINPUT34), .ZN(n412) );
  NAND2_X1 U539 ( .A1(n464), .A2(n465), .ZN(n463) );
  AND2_X2 U540 ( .A1(n425), .A2(n423), .ZN(n422) );
  NAND2_X1 U541 ( .A1(n424), .A2(KEYINPUT45), .ZN(n423) );
  NAND2_X1 U542 ( .A1(n426), .A2(n580), .ZN(n424) );
  NAND2_X1 U543 ( .A1(n593), .A2(n357), .ZN(n426) );
  NAND2_X1 U544 ( .A1(n589), .A2(KEYINPUT44), .ZN(n428) );
  INV_X1 U545 ( .A(n430), .ZN(n573) );
  NAND2_X1 U546 ( .A1(n430), .A2(n566), .ZN(n451) );
  NAND2_X1 U547 ( .A1(n351), .A2(n607), .ZN(n576) );
  AND2_X1 U548 ( .A1(n431), .A2(n639), .ZN(n434) );
  XNOR2_X2 U549 ( .A(n554), .B(G472), .ZN(n612) );
  NAND2_X1 U550 ( .A1(n603), .A2(n442), .ZN(n441) );
  XNOR2_X2 U551 ( .A(n460), .B(n523), .ZN(n603) );
  INV_X1 U552 ( .A(n603), .ZN(n439) );
  NAND2_X1 U553 ( .A1(n715), .A2(n642), .ZN(n460) );
  NAND2_X1 U554 ( .A1(n758), .A2(n472), .ZN(n470) );
  NAND2_X1 U555 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U556 ( .A(n609), .B(n443), .ZN(n619) );
  NAND2_X1 U557 ( .A1(n770), .A2(n769), .ZN(n444) );
  XNOR2_X1 U558 ( .A(n766), .B(n586), .ZN(n591) );
  NAND2_X1 U559 ( .A1(n445), .A2(n627), .ZN(n637) );
  NAND2_X1 U560 ( .A1(n625), .A2(n468), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n446), .B(n504), .ZN(n507) );
  XNOR2_X1 U562 ( .A(n503), .B(n356), .ZN(n446) );
  XNOR2_X1 U563 ( .A(n638), .B(KEYINPUT72), .ZN(n464) );
  INV_X1 U564 ( .A(n758), .ZN(n454) );
  NOR2_X2 U565 ( .A1(n585), .A2(n567), .ZN(n583) );
  AND2_X1 U566 ( .A1(n376), .A2(n759), .ZN(n748) );
  INV_X1 U567 ( .A(KEYINPUT45), .ZN(n456) );
  OR2_X2 U568 ( .A1(n768), .A2(n457), .ZN(n458) );
  NAND2_X1 U569 ( .A1(n458), .A2(KEYINPUT66), .ZN(n588) );
  NAND2_X1 U570 ( .A1(n375), .A2(G472), .ZN(n644) );
  NAND2_X1 U571 ( .A1(n379), .A2(G210), .ZN(n717) );
  NAND2_X1 U572 ( .A1(n375), .A2(G475), .ZN(n729) );
  NAND2_X1 U573 ( .A1(n462), .A2(G217), .ZN(n739) );
  NAND2_X1 U574 ( .A1(n379), .A2(G478), .ZN(n733) );
  NAND2_X1 U575 ( .A1(n462), .A2(G469), .ZN(n724) );
  INV_X1 U576 ( .A(n465), .ZN(n709) );
  NAND2_X1 U577 ( .A1(n468), .A2(n706), .ZN(n697) );
  NAND2_X1 U578 ( .A1(n468), .A2(n703), .ZN(n701) );
  NAND2_X1 U579 ( .A1(n470), .A2(n471), .ZN(n469) );
  INV_X1 U580 ( .A(KEYINPUT2), .ZN(n472) );
  XNOR2_X2 U581 ( .A(n474), .B(n549), .ZN(n653) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U583 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U584 ( .A(n739), .B(n738), .ZN(n741) );
  NOR2_X2 U585 ( .A1(n624), .A2(n532), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n564), .A2(n651), .ZN(n572) );
  NOR2_X1 U587 ( .A1(n572), .A2(n598), .ZN(n555) );
  XNOR2_X1 U588 ( .A(n384), .B(n714), .ZN(n716) );
  AND2_X1 U589 ( .A1(G227), .A2(n759), .ZN(n475) );
  INV_X1 U590 ( .A(KEYINPUT48), .ZN(n641) );
  XNOR2_X1 U591 ( .A(n486), .B(n513), .ZN(n487) );
  XNOR2_X1 U592 ( .A(n537), .B(n487), .ZN(n553) );
  XNOR2_X1 U593 ( .A(n513), .B(n355), .ZN(n514) );
  INV_X1 U594 ( .A(n650), .ZN(n640) );
  INV_X1 U595 ( .A(KEYINPUT122), .ZN(n686) );
  XNOR2_X1 U596 ( .A(n688), .B(n687), .ZN(G75) );
  XNOR2_X2 U597 ( .A(G143), .B(KEYINPUT64), .ZN(n476) );
  XNOR2_X2 U598 ( .A(n476), .B(G128), .ZN(n498) );
  NOR2_X2 U599 ( .A1(G953), .A2(G237), .ZN(n505) );
  NAND2_X1 U600 ( .A1(n505), .A2(G210), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U602 ( .A(n481), .B(KEYINPUT75), .Z(n483) );
  XNOR2_X1 U603 ( .A(n483), .B(n482), .ZN(n486) );
  XOR2_X1 U604 ( .A(G113), .B(G116), .Z(n485) );
  XNOR2_X1 U605 ( .A(G119), .B(KEYINPUT3), .ZN(n484) );
  XNOR2_X1 U606 ( .A(n485), .B(n484), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U609 ( .A(n493), .B(n492), .Z(n496) );
  NAND2_X1 U610 ( .A1(G234), .A2(n759), .ZN(n494) );
  NAND2_X1 U611 ( .A1(G217), .A2(n545), .ZN(n495) );
  XNOR2_X1 U612 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U613 ( .A(n377), .B(n497), .ZN(n734) );
  NOR2_X1 U614 ( .A1(G902), .A2(n734), .ZN(n500) );
  XNOR2_X1 U615 ( .A(KEYINPUT107), .B(G478), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n571) );
  XOR2_X1 U617 ( .A(G131), .B(G122), .Z(n502) );
  XNOR2_X1 U618 ( .A(G104), .B(G113), .ZN(n501) );
  XNOR2_X1 U619 ( .A(n502), .B(n501), .ZN(n504) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n503) );
  NAND2_X1 U621 ( .A1(n505), .A2(G214), .ZN(n506) );
  XNOR2_X1 U622 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U623 ( .A(n754), .B(n508), .ZN(n726) );
  NOR2_X1 U624 ( .A1(G902), .A2(n726), .ZN(n509) );
  NAND2_X1 U625 ( .A1(n571), .A2(n569), .ZN(n630) );
  XOR2_X1 U626 ( .A(n630), .B(KEYINPUT76), .Z(n557) );
  XOR2_X1 U627 ( .A(KEYINPUT90), .B(G107), .Z(n511) );
  XNOR2_X1 U628 ( .A(G104), .B(G101), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U630 ( .A1(G224), .A2(n759), .ZN(n517) );
  XOR2_X1 U631 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n521) );
  NAND2_X1 U632 ( .A1(G210), .A2(n524), .ZN(n520) );
  XNOR2_X1 U633 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U634 ( .A(KEYINPUT77), .B(n522), .Z(n523) );
  NAND2_X1 U635 ( .A1(n524), .A2(G214), .ZN(n525) );
  XOR2_X1 U636 ( .A(KEYINPUT94), .B(n525), .Z(n665) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n527) );
  XNOR2_X1 U638 ( .A(n527), .B(n526), .ZN(n529) );
  NAND2_X1 U639 ( .A1(n529), .A2(G952), .ZN(n528) );
  XOR2_X1 U640 ( .A(KEYINPUT96), .B(n528), .Z(n679) );
  NAND2_X1 U641 ( .A1(n759), .A2(n679), .ZN(n597) );
  INV_X1 U642 ( .A(n597), .ZN(n531) );
  XNOR2_X1 U643 ( .A(G898), .B(KEYINPUT97), .ZN(n747) );
  NAND2_X1 U644 ( .A1(G953), .A2(n747), .ZN(n744) );
  NAND2_X1 U645 ( .A1(G902), .A2(n529), .ZN(n594) );
  NOR2_X1 U646 ( .A1(n744), .A2(n594), .ZN(n530) );
  NOR2_X1 U647 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U648 ( .A(KEYINPUT98), .B(n540), .ZN(n756) );
  XNOR2_X1 U649 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U650 ( .A(KEYINPUT71), .B(G469), .ZN(n538) );
  XNOR2_X2 U651 ( .A(n539), .B(n538), .ZN(n615) );
  XOR2_X1 U652 ( .A(KEYINPUT24), .B(G128), .Z(n542) );
  XNOR2_X1 U653 ( .A(G110), .B(G119), .ZN(n541) );
  XNOR2_X1 U654 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U655 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n548) );
  NAND2_X1 U656 ( .A1(G234), .A2(n642), .ZN(n546) );
  XNOR2_X1 U657 ( .A(KEYINPUT20), .B(n546), .ZN(n550) );
  NAND2_X1 U658 ( .A1(n550), .A2(G217), .ZN(n547) );
  XNOR2_X1 U659 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U660 ( .A1(n550), .A2(G221), .ZN(n551) );
  XNOR2_X1 U661 ( .A(n551), .B(KEYINPUT102), .ZN(n552) );
  XNOR2_X1 U662 ( .A(KEYINPUT21), .B(n552), .ZN(n654) );
  NOR2_X1 U663 ( .A1(G902), .A2(n553), .ZN(n554) );
  XNOR2_X1 U664 ( .A(n555), .B(KEYINPUT33), .ZN(n673) );
  NOR2_X2 U665 ( .A1(n573), .A2(n673), .ZN(n556) );
  XNOR2_X1 U666 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n558) );
  XNOR2_X2 U667 ( .A(n559), .B(n558), .ZN(n766) );
  NAND2_X1 U668 ( .A1(n766), .A2(KEYINPUT85), .ZN(n560) );
  NAND2_X1 U669 ( .A1(n560), .A2(KEYINPUT44), .ZN(n563) );
  INV_X1 U670 ( .A(KEYINPUT85), .ZN(n561) );
  NAND2_X1 U671 ( .A1(n561), .A2(KEYINPUT66), .ZN(n562) );
  NAND2_X1 U672 ( .A1(n563), .A2(n562), .ZN(n580) );
  INV_X1 U673 ( .A(n654), .ZN(n565) );
  NOR2_X1 U674 ( .A1(n571), .A2(n569), .ZN(n667) );
  AND2_X1 U675 ( .A1(n565), .A2(n667), .ZN(n566) );
  INV_X1 U676 ( .A(n598), .ZN(n567) );
  XNOR2_X1 U677 ( .A(n583), .B(KEYINPUT84), .ZN(n568) );
  INV_X1 U678 ( .A(n653), .ZN(n581) );
  INV_X1 U679 ( .A(n569), .ZN(n570) );
  NOR2_X1 U680 ( .A1(n571), .A2(n570), .ZN(n618) );
  AND2_X1 U681 ( .A1(n571), .A2(n570), .ZN(n706) );
  NOR2_X1 U682 ( .A1(n618), .A2(n706), .ZN(n628) );
  OR2_X1 U683 ( .A1(n612), .A2(n572), .ZN(n661) );
  NOR2_X1 U684 ( .A1(n573), .A2(n661), .ZN(n574) );
  XOR2_X1 U685 ( .A(KEYINPUT31), .B(n574), .Z(n707) );
  INV_X1 U686 ( .A(n612), .ZN(n656) );
  NAND2_X1 U687 ( .A1(n651), .A2(n615), .ZN(n575) );
  NOR2_X1 U688 ( .A1(n656), .A2(n576), .ZN(n692) );
  NOR2_X1 U689 ( .A1(n707), .A2(n692), .ZN(n577) );
  NOR2_X1 U690 ( .A1(n628), .A2(n577), .ZN(n578) );
  NOR2_X1 U691 ( .A1(n689), .A2(n578), .ZN(n579) );
  NOR2_X1 U692 ( .A1(n640), .A2(n581), .ZN(n582) );
  INV_X1 U693 ( .A(KEYINPUT67), .ZN(n586) );
  OR2_X1 U694 ( .A1(n766), .A2(KEYINPUT85), .ZN(n587) );
  NAND2_X1 U695 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U696 ( .A(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U697 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U698 ( .A1(n592), .A2(KEYINPUT66), .ZN(n593) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT109), .ZN(n690) );
  NOR2_X1 U700 ( .A1(G900), .A2(n594), .ZN(n595) );
  NAND2_X1 U701 ( .A1(G953), .A2(n595), .ZN(n596) );
  NAND2_X1 U702 ( .A1(n597), .A2(n596), .ZN(n605) );
  NOR2_X1 U703 ( .A1(n665), .A2(n650), .ZN(n600) );
  NAND2_X1 U704 ( .A1(n639), .A2(n600), .ZN(n601) );
  XNOR2_X1 U705 ( .A(KEYINPUT43), .B(n601), .ZN(n602) );
  XOR2_X1 U706 ( .A(KEYINPUT111), .B(n602), .Z(n604) );
  OR2_X1 U707 ( .A1(n612), .A2(n665), .ZN(n606) );
  XOR2_X1 U708 ( .A(KEYINPUT38), .B(KEYINPUT74), .Z(n608) );
  XNOR2_X1 U709 ( .A(n631), .B(n608), .ZN(n664) );
  AND2_X1 U710 ( .A1(n619), .A2(n706), .ZN(n712) );
  NOR2_X1 U711 ( .A1(n665), .A2(n664), .ZN(n670) );
  NAND2_X1 U712 ( .A1(n670), .A2(n667), .ZN(n611) );
  XOR2_X1 U713 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n610) );
  XNOR2_X1 U714 ( .A(n611), .B(n610), .ZN(n683) );
  XNOR2_X1 U715 ( .A(KEYINPUT28), .B(n614), .ZN(n616) );
  NAND2_X1 U716 ( .A1(n616), .A2(n615), .ZN(n623) );
  NOR2_X1 U717 ( .A1(n683), .A2(n623), .ZN(n617) );
  XOR2_X1 U718 ( .A(KEYINPUT42), .B(n617), .Z(n769) );
  XNOR2_X1 U719 ( .A(n620), .B(KEYINPUT40), .ZN(n770) );
  XOR2_X1 U720 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n621) );
  INV_X1 U721 ( .A(n628), .ZN(n669) );
  NAND2_X1 U722 ( .A1(n621), .A2(n669), .ZN(n622) );
  XNOR2_X1 U723 ( .A(n622), .B(KEYINPUT73), .ZN(n625) );
  NAND2_X1 U724 ( .A1(n626), .A2(KEYINPUT47), .ZN(n627) );
  INV_X1 U725 ( .A(KEYINPUT79), .ZN(n635) );
  NAND2_X1 U726 ( .A1(KEYINPUT47), .A2(n628), .ZN(n633) );
  NOR2_X1 U727 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U728 ( .A1(n633), .A2(n700), .ZN(n634) );
  XNOR2_X1 U729 ( .A(n634), .B(n635), .ZN(n636) );
  NOR2_X1 U730 ( .A1(G952), .A2(n759), .ZN(n646) );
  INV_X1 U731 ( .A(n736), .ZN(n740) );
  XNOR2_X1 U732 ( .A(KEYINPUT87), .B(KEYINPUT115), .ZN(n647) );
  XNOR2_X1 U733 ( .A(n647), .B(KEYINPUT63), .ZN(n648) );
  XNOR2_X1 U734 ( .A(n649), .B(n648), .ZN(G57) );
  NOR2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U736 ( .A(KEYINPUT50), .B(n652), .Z(n659) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n655), .B(KEYINPUT49), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT51), .B(n662), .ZN(n663) );
  NOR2_X1 U743 ( .A1(n683), .A2(n663), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(KEYINPUT121), .ZN(n672) );
  AND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n674) );
  NOR2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT52), .B(n677), .Z(n678) );
  NAND2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n683), .A2(n673), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n686), .B(KEYINPUT53), .ZN(n687) );
  XOR2_X1 U755 ( .A(n689), .B(G101), .Z(G3) );
  INV_X1 U756 ( .A(n690), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n692), .A2(n703), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(G104), .ZN(G6) );
  XOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U760 ( .A1(n692), .A2(n706), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(G107), .B(n695), .ZN(G9) );
  XOR2_X1 U763 ( .A(G110), .B(n696), .Z(G12) );
  XOR2_X1 U764 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U766 ( .A(G128), .B(n699), .ZN(G30) );
  XNOR2_X1 U767 ( .A(G143), .B(n700), .ZN(G45) );
  XOR2_X1 U768 ( .A(G146), .B(KEYINPUT117), .Z(n702) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(G48) );
  NAND2_X1 U770 ( .A1(n707), .A2(n703), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n704), .B(KEYINPUT118), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G113), .B(n705), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(G116), .ZN(G18) );
  XOR2_X1 U775 ( .A(KEYINPUT119), .B(KEYINPUT37), .Z(n711) );
  XNOR2_X1 U776 ( .A(G125), .B(n709), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n711), .B(n710), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(n712), .Z(n713) );
  XNOR2_X1 U779 ( .A(KEYINPUT120), .B(n713), .ZN(G36) );
  XOR2_X1 U780 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n714) );
  XNOR2_X1 U781 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n718), .A2(n740), .ZN(n720) );
  XNOR2_X1 U783 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n719) );
  XNOR2_X1 U784 ( .A(n720), .B(n719), .ZN(G51) );
  XOR2_X1 U785 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n722) );
  NOR2_X1 U786 ( .A1(n736), .A2(n725), .ZN(G54) );
  XNOR2_X1 U787 ( .A(n726), .B(KEYINPUT88), .ZN(n727) );
  XNOR2_X1 U788 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U789 ( .A1(n730), .A2(n740), .ZN(n732) );
  XOR2_X1 U790 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n731) );
  XNOR2_X1 U791 ( .A(n732), .B(n731), .ZN(G60) );
  XNOR2_X1 U792 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(G63) );
  INV_X1 U794 ( .A(n737), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n751) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n745) );
  XOR2_X1 U798 ( .A(KEYINPUT61), .B(n745), .Z(n746) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n749) );
  NOR2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U802 ( .A(KEYINPUT126), .B(n752), .ZN(G69) );
  XOR2_X1 U803 ( .A(n754), .B(n753), .Z(n755) );
  XOR2_X1 U804 ( .A(n756), .B(n755), .Z(n761) );
  XOR2_X1 U805 ( .A(KEYINPUT127), .B(n761), .Z(n757) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U808 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n765), .A2(n764), .ZN(G72) );
  XNOR2_X1 U812 ( .A(n352), .B(G122), .ZN(G24) );
  XNOR2_X1 U813 ( .A(G140), .B(n767), .ZN(G42) );
  XOR2_X1 U814 ( .A(n768), .B(G119), .Z(G21) );
  XNOR2_X1 U815 ( .A(G137), .B(n769), .ZN(G39) );
  XNOR2_X1 U816 ( .A(G131), .B(n770), .ZN(G33) );
endmodule

