

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580;

  INV_X1 U319 ( .A(KEYINPUT55), .ZN(n467) );
  XNOR2_X1 U320 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U321 ( .A(n392), .B(n349), .ZN(n350) );
  XNOR2_X1 U322 ( .A(n452), .B(KEYINPUT109), .ZN(n453) );
  XNOR2_X1 U323 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U324 ( .A(G92GAT), .ZN(n431) );
  XNOR2_X1 U325 ( .A(n454), .B(n453), .ZN(n460) );
  XNOR2_X1 U326 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U327 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n405) );
  XNOR2_X1 U328 ( .A(n434), .B(n433), .ZN(n442) );
  XNOR2_X1 U329 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U330 ( .A(n406), .B(n405), .ZN(n508) );
  XNOR2_X1 U331 ( .A(n473), .B(G190GAT), .ZN(n474) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XNOR2_X1 U334 ( .A(n446), .B(n445), .ZN(G1330GAT) );
  XNOR2_X1 U335 ( .A(G57GAT), .B(G64GAT), .ZN(n287) );
  XNOR2_X1 U336 ( .A(n287), .B(KEYINPUT13), .ZN(n427) );
  XOR2_X1 U337 ( .A(n427), .B(G211GAT), .Z(n289) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G71GAT), .Z(n352) );
  XNOR2_X1 U339 ( .A(n352), .B(G155GAT), .ZN(n288) );
  XNOR2_X1 U340 ( .A(n289), .B(n288), .ZN(n295) );
  XOR2_X1 U341 ( .A(KEYINPUT68), .B(G8GAT), .Z(n291) );
  XNOR2_X1 U342 ( .A(G22GAT), .B(G1GAT), .ZN(n290) );
  XNOR2_X1 U343 ( .A(n291), .B(n290), .ZN(n422) );
  XOR2_X1 U344 ( .A(n422), .B(KEYINPUT12), .Z(n293) );
  NAND2_X1 U345 ( .A1(G231GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U347 ( .A(n295), .B(n294), .Z(n303) );
  XOR2_X1 U348 ( .A(KEYINPUT79), .B(G78GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(G183GAT), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n299) );
  XNOR2_X1 U352 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n573) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n304), .B(KEYINPUT86), .ZN(n305) );
  XOR2_X1 U358 ( .A(n305), .B(KEYINPUT3), .Z(n307) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(G148GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n335) );
  XOR2_X1 U361 ( .A(KEYINPUT1), .B(G57GAT), .Z(n309) );
  XNOR2_X1 U362 ( .A(G134GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n314) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(KEYINPUT75), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n310), .B(G85GAT), .ZN(n401) );
  XOR2_X1 U366 ( .A(n401), .B(KEYINPUT5), .Z(n312) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n314), .B(n313), .Z(n321) );
  XNOR2_X1 U370 ( .A(G120GAT), .B(G127GAT), .ZN(n316) );
  XOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .Z(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n351) );
  XOR2_X1 U373 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n318) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n351), .B(n319), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n335), .B(n322), .ZN(n379) );
  XOR2_X1 U379 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n324) );
  XNOR2_X1 U380 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n339) );
  XOR2_X1 U382 ( .A(G204GAT), .B(G78GAT), .Z(n430) );
  XOR2_X1 U383 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n326) );
  XNOR2_X1 U384 ( .A(G22GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n430), .B(n327), .ZN(n329) );
  AND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n332) );
  XOR2_X1 U389 ( .A(G211GAT), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U390 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n363) );
  XOR2_X1 U392 ( .A(n332), .B(n363), .Z(n337) );
  XOR2_X1 U393 ( .A(G162GAT), .B(KEYINPUT72), .Z(n334) );
  XNOR2_X1 U394 ( .A(G50GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n395) );
  XNOR2_X1 U396 ( .A(n335), .B(n395), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U398 ( .A(n339), .B(n338), .Z(n370) );
  BUF_X1 U399 ( .A(n370), .Z(n466) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n340), .B(KEYINPUT19), .ZN(n341) );
  XOR2_X1 U402 ( .A(n341), .B(KEYINPUT17), .Z(n343) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(G176GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n364) );
  XOR2_X1 U405 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n345) );
  XNOR2_X1 U406 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n364), .B(n346), .Z(n348) );
  XNOR2_X1 U409 ( .A(G190GAT), .B(G99GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n355) );
  XOR2_X1 U411 ( .A(G43GAT), .B(G134GAT), .Z(n392) );
  AND2_X1 U412 ( .A1(G227GAT), .A2(G233GAT), .ZN(n349) );
  XOR2_X1 U413 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n369) );
  INV_X1 U415 ( .A(n369), .ZN(n472) );
  INV_X1 U416 ( .A(n472), .ZN(n524) );
  XNOR2_X1 U417 ( .A(G36GAT), .B(G190GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(G92GAT), .ZN(n400) );
  XOR2_X1 U419 ( .A(G64GAT), .B(n400), .Z(n358) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(G204GAT), .Z(n360) );
  XNOR2_X1 U423 ( .A(G8GAT), .B(G218GAT), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U425 ( .A(n362), .B(n361), .Z(n366) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n462) );
  INV_X1 U428 ( .A(n462), .ZN(n512) );
  NAND2_X1 U429 ( .A1(n524), .A2(n512), .ZN(n367) );
  NAND2_X1 U430 ( .A1(n466), .A2(n367), .ZN(n368) );
  XNOR2_X1 U431 ( .A(KEYINPUT25), .B(n368), .ZN(n376) );
  NOR2_X1 U432 ( .A1(n370), .A2(n369), .ZN(n372) );
  XNOR2_X1 U433 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U435 ( .A(KEYINPUT94), .B(n373), .Z(n564) );
  XOR2_X1 U436 ( .A(n462), .B(KEYINPUT27), .Z(n380) );
  NAND2_X1 U437 ( .A1(n564), .A2(n380), .ZN(n374) );
  XOR2_X1 U438 ( .A(KEYINPUT96), .B(n374), .Z(n375) );
  NOR2_X1 U439 ( .A1(n376), .A2(n375), .ZN(n377) );
  XOR2_X1 U440 ( .A(n377), .B(KEYINPUT97), .Z(n378) );
  NOR2_X1 U441 ( .A1(n379), .A2(n378), .ZN(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT90), .B(n379), .ZN(n510) );
  NAND2_X1 U443 ( .A1(n380), .A2(n510), .ZN(n381) );
  XOR2_X1 U444 ( .A(KEYINPUT92), .B(n381), .Z(n538) );
  XNOR2_X1 U445 ( .A(n466), .B(KEYINPUT28), .ZN(n486) );
  NAND2_X1 U446 ( .A1(n538), .A2(n486), .ZN(n522) );
  XNOR2_X1 U447 ( .A(KEYINPUT83), .B(n472), .ZN(n382) );
  NOR2_X1 U448 ( .A1(n522), .A2(n382), .ZN(n383) );
  XOR2_X1 U449 ( .A(KEYINPUT93), .B(n383), .Z(n384) );
  NOR2_X2 U450 ( .A1(n385), .A2(n384), .ZN(n479) );
  NOR2_X1 U451 ( .A1(n573), .A2(n479), .ZN(n387) );
  INV_X1 U452 ( .A(KEYINPUT99), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n404) );
  XOR2_X1 U454 ( .A(G99GAT), .B(G106GAT), .Z(n426) );
  XOR2_X1 U455 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n389) );
  XNOR2_X1 U456 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U458 ( .A(n426), .B(n390), .Z(n394) );
  XNOR2_X1 U459 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n391), .B(KEYINPUT7), .ZN(n423) );
  XNOR2_X1 U461 ( .A(n423), .B(n392), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U463 ( .A(n395), .B(KEYINPUT74), .Z(n397) );
  NAND2_X1 U464 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n403) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n549) );
  XNOR2_X1 U469 ( .A(n549), .B(KEYINPUT76), .ZN(n533) );
  XNOR2_X1 U470 ( .A(KEYINPUT36), .B(n533), .ZN(n576) );
  NAND2_X1 U471 ( .A1(n404), .A2(n576), .ZN(n406) );
  XOR2_X1 U472 ( .A(G36GAT), .B(G29GAT), .Z(n408) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(G43GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U475 ( .A(G15GAT), .B(G197GAT), .Z(n410) );
  XNOR2_X1 U476 ( .A(G169GAT), .B(G141GAT), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U479 ( .A(KEYINPUT66), .B(KEYINPUT70), .Z(n414) );
  NAND2_X1 U480 ( .A1(G229GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U482 ( .A(KEYINPUT69), .B(n415), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U484 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n419) );
  XNOR2_X1 U485 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U487 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n497) );
  XOR2_X1 U490 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n430), .B(G85GAT), .ZN(n432) );
  XOR2_X1 U494 ( .A(G148GAT), .B(G120GAT), .Z(n436) );
  XNOR2_X1 U495 ( .A(G176GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n438) );
  XNOR2_X1 U498 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n570) );
  NOR2_X1 U502 ( .A1(n497), .A2(n570), .ZN(n480) );
  NAND2_X1 U503 ( .A1(n508), .A2(n480), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n443), .B(KEYINPUT38), .ZN(n444) );
  XNOR2_X1 U505 ( .A(KEYINPUT101), .B(n444), .ZN(n494) );
  NAND2_X1 U506 ( .A1(n494), .A2(n524), .ZN(n446) );
  INV_X1 U507 ( .A(KEYINPUT108), .ZN(n450) );
  XNOR2_X1 U508 ( .A(KEYINPUT41), .B(n570), .ZN(n496) );
  NOR2_X1 U509 ( .A1(n497), .A2(n496), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n447), .B(KEYINPUT46), .ZN(n448) );
  NOR2_X1 U511 ( .A1(n448), .A2(n573), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U513 ( .A1(n549), .A2(n451), .ZN(n454) );
  INV_X1 U514 ( .A(KEYINPUT47), .ZN(n452) );
  XOR2_X1 U515 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n456) );
  NAND2_X1 U516 ( .A1(n573), .A2(n576), .ZN(n455) );
  XOR2_X1 U517 ( .A(n456), .B(n455), .Z(n457) );
  NOR2_X1 U518 ( .A1(n570), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n458), .A2(n497), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT48), .B(n461), .Z(n540) );
  NOR2_X1 U522 ( .A1(n540), .A2(n462), .ZN(n464) );
  INV_X1 U523 ( .A(KEYINPUT54), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n510), .A2(n465), .ZN(n563) );
  NAND2_X1 U526 ( .A1(n563), .A2(n466), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n468) );
  NOR2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n561) );
  NAND2_X1 U529 ( .A1(n561), .A2(n533), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n473) );
  INV_X1 U531 ( .A(n573), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n476), .A2(n533), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n498) );
  AND2_X1 U535 ( .A1(n480), .A2(n498), .ZN(n487) );
  NAND2_X1 U536 ( .A1(n487), .A2(n510), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n512), .A2(n487), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U542 ( .A1(n487), .A2(n524), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n486), .ZN(n516) );
  NAND2_X1 U545 ( .A1(n487), .A2(n516), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT98), .B(KEYINPUT102), .Z(n490) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n510), .A2(n494), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n494), .A2(n512), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n494), .A2(n516), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U556 ( .A(n497), .ZN(n566) );
  NOR2_X1 U557 ( .A1(n496), .A2(n566), .ZN(n509) );
  AND2_X1 U558 ( .A1(n509), .A2(n498), .ZN(n504) );
  NAND2_X1 U559 ( .A1(n510), .A2(n504), .ZN(n499) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(n499), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  XOR2_X1 U562 ( .A(G64GAT), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U563 ( .A1(n504), .A2(n512), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n524), .A2(n504), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U568 ( .A1(n504), .A2(n516), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G78GAT), .B(n507), .ZN(G1335GAT) );
  AND2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  XOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U575 ( .A1(n517), .A2(n512), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1337GAT) );
  NAND2_X1 U577 ( .A1(n524), .A2(n517), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(KEYINPUT106), .ZN(n521) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U584 ( .A1(n540), .A2(n522), .ZN(n523) );
  NAND2_X1 U585 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n525), .Z(n534) );
  NAND2_X1 U587 ( .A1(n534), .A2(n566), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n528) );
  INV_X1 U590 ( .A(n496), .ZN(n558) );
  NAND2_X1 U591 ( .A1(n534), .A2(n558), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U593 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n531) );
  NAND2_X1 U595 ( .A1(n573), .A2(n534), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(G134GAT), .B(n537), .Z(G1343GAT) );
  NAND2_X1 U602 ( .A1(n564), .A2(n538), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n566), .A2(n550), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 U606 ( .A1(n558), .A2(n550), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT114), .Z(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n573), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U615 ( .A(G162GAT), .B(KEYINPUT117), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1347GAT) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n561), .A2(n566), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n573), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(n565), .Z(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n575), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1355GAT) );
endmodule

