//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(G160));
  NAND2_X1  g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n471), .A2(new_n474), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n492), .B(new_n493), .C1(new_n473), .C2(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n463), .B2(new_n492), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n463), .A2(new_n503), .A3(G126), .A4(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n508), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(G62), .B1(new_n510), .B2(new_n508), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n509), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n518), .B1(new_n527), .B2(G651), .ZN(G166));
  NAND3_X1  g103(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT71), .Z(new_n530));
  INV_X1    g105(.A(new_n513), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(new_n511), .B1(new_n523), .B2(new_n509), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n522), .B1(new_n531), .B2(new_n511), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n530), .A2(new_n538), .ZN(G168));
  XOR2_X1   g114(.A(KEYINPUT72), .B(G52), .Z(new_n540));
  AOI22_X1  g115(.A1(new_n532), .A2(G90), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT73), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n544), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n514), .A2(new_n550), .B1(new_n516), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT74), .Z(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n524), .B(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n516), .A2(KEYINPUT9), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n516), .B2(new_n566), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(new_n568), .B1(G91), .B2(new_n532), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n516), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n532), .A2(G87), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G288));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n523), .B2(new_n509), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n514), .A2(new_n585), .B1(new_n586), .B2(new_n516), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n532), .A2(G85), .B1(new_n534), .B2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n544), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT76), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n532), .A2(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n534), .A2(G54), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n561), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n561), .A2(new_n602), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n544), .B1(new_n608), .B2(new_n604), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n598), .A2(new_n599), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT77), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n595), .B1(new_n612), .B2(new_n594), .ZN(G284));
  AOI21_X1  g188(.A(new_n595), .B1(new_n612), .B2(new_n594), .ZN(G321));
  OR3_X1    g189(.A1(G168), .A2(KEYINPUT78), .A3(new_n594), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(G168), .B2(new_n594), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n565), .A2(new_n569), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n617), .ZN(G297));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n483), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n631));
  OR3_X1    g206(.A1(new_n631), .A2(new_n464), .A3(G111), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n464), .B2(G111), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n630), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n471), .A2(new_n474), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n461), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n637), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n670), .B(KEYINPUT17), .Z(new_n675));
  OAI211_X1 g250(.A(new_n672), .B(new_n674), .C1(new_n669), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n668), .A3(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n669), .A3(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n684), .A2(new_n689), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n692));
  AOI211_X1 g267(.A(new_n688), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G19), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n553), .B2(new_n702), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1341), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n702), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(G1966), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n636), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT96), .B(KEYINPUT31), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G11), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(G28), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT98), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n718), .A2(KEYINPUT98), .B1(new_n716), .B2(G28), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n712), .A2(new_n713), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n709), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n709), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT29), .B(G2090), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2078), .ZN(new_n727));
  NOR2_X1   g302(.A1(G164), .A2(new_n709), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G27), .B2(new_n709), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n722), .B(new_n726), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n708), .B(new_n730), .C1(G1966), .C2(new_n707), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n709), .A2(G26), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  OR2_X1    g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  INV_X1    g311(.A(G128), .ZN(new_n737));
  INV_X1    g312(.A(G140), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n737), .A2(new_n480), .B1(new_n465), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n741), .A2(KEYINPUT92), .A3(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT92), .B1(new_n741), .B2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n733), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n747), .B2(KEYINPUT24), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(KEYINPUT24), .B2(new_n747), .ZN(new_n749));
  INV_X1    g324(.A(G160), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n709), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n702), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT100), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n617), .B2(new_n702), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT101), .B(G1956), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n760), .B(new_n761), .C1(new_n727), .C2(new_n729), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n731), .A2(new_n746), .A3(new_n753), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n612), .B2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT90), .B(G1348), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n709), .A2(G32), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n483), .A2(G141), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  INV_X1    g347(.A(G129), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n480), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n461), .A2(G105), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n770), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n709), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT95), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT27), .ZN(new_n779));
  INV_X1    g354(.A(G1996), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n763), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n588), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g360(.A(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n702), .A2(G23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n577), .B2(new_n702), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G22), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G166), .B2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n791), .B1(G1971), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n787), .B(new_n794), .C1(G1971), .C2(new_n793), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n797));
  OR2_X1    g372(.A1(G16), .A2(G24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G290), .B2(new_n702), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1986), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n803));
  INV_X1    g378(.A(G131), .ZN(new_n804));
  INV_X1    g379(.A(G119), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(new_n465), .B2(new_n804), .C1(new_n805), .C2(new_n480), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  AOI211_X1 g386(.A(KEYINPUT89), .B(new_n810), .C1(new_n799), .C2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n796), .A2(new_n797), .A3(new_n801), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n638), .A2(G127), .ZN(new_n816));
  INV_X1    g391(.A(G115), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n460), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT93), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n464), .B1(new_n818), .B2(KEYINPUT93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n483), .A2(G139), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G29), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G29), .B2(G33), .ZN(new_n829));
  INV_X1    g404(.A(G2072), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT94), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n702), .A2(G5), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G171), .B2(new_n702), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT99), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n835), .A2(G1961), .B1(new_n752), .B2(new_n751), .ZN(new_n836));
  OAI221_X1 g411(.A(new_n836), .B1(G1961), .B2(new_n835), .C1(new_n830), .C2(new_n829), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n813), .A2(new_n814), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n782), .A2(new_n815), .A3(new_n838), .A4(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  AOI22_X1  g416(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n544), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n514), .A2(new_n844), .B1(new_n516), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n553), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n612), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n620), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT103), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n849), .B(new_n553), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n862), .A3(KEYINPUT39), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT104), .B(G860), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n847), .A2(new_n867), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n776), .B1(new_n827), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n821), .A2(new_n826), .ZN(new_n875));
  INV_X1    g450(.A(new_n776), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(KEYINPUT106), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n874), .A2(new_n740), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n740), .B1(new_n874), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(G164), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n741), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n874), .A2(new_n740), .A3(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n506), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n806), .B(KEYINPUT107), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n640), .ZN(new_n887));
  OR2_X1    g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n889));
  INV_X1    g464(.A(G142), .ZN(new_n890));
  INV_X1    g465(.A(G130), .ZN(new_n891));
  OAI221_X1 g466(.A(new_n889), .B1(new_n465), .B2(new_n890), .C1(new_n891), .C2(new_n480), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n893), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n636), .B(new_n487), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT105), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G160), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n880), .A2(new_n884), .A3(new_n898), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n900), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n872), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n904), .ZN(new_n910));
  INV_X1    g485(.A(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n906), .A4(new_n905), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n909), .A2(new_n913), .ZN(G395));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n851), .A2(new_n620), .A3(new_n612), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n622), .A2(new_n861), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n600), .A2(new_n606), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G299), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n617), .A2(new_n606), .A3(new_n600), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT109), .B1(new_n922), .B2(KEYINPUT41), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n919), .A2(G299), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n600), .A2(new_n606), .B1(new_n565), .B2(new_n569), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT41), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n921), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n925), .B1(new_n931), .B2(KEYINPUT109), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n924), .B(KEYINPUT110), .C1(new_n932), .C2(new_n918), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  INV_X1    g509(.A(new_n918), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n928), .B2(new_n930), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n935), .B(new_n936), .C1(new_n938), .C2(new_n925), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n933), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n933), .B2(new_n939), .ZN(new_n941));
  XNOR2_X1  g516(.A(G290), .B(G303), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n577), .B(KEYINPUT111), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(G305), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n942), .A2(new_n944), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n940), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n941), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G868), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n915), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n594), .B1(new_n843), .B2(new_n846), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n594), .B1(new_n941), .B2(new_n951), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n941), .A2(new_n951), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT113), .B(new_n957), .C1(new_n958), .C2(new_n940), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(G295));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(G331));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  XNOR2_X1  g537(.A(G301), .B(G286), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n861), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(G301), .B(G168), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n851), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n938), .B2(new_n925), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n964), .A2(new_n966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n923), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n970), .A3(new_n948), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n970), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n946), .A2(new_n947), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n967), .A2(new_n931), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n967), .A2(new_n922), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n971), .A3(new_n906), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n962), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n971), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n973), .A2(new_n906), .A3(new_n980), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n988), .B2(new_n962), .ZN(G397));
  NAND2_X1  g564(.A1(new_n477), .A2(G2105), .ZN(new_n990));
  INV_X1    g565(.A(new_n467), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT114), .B(G40), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n478), .A2(KEYINPUT115), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n506), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n740), .A2(new_n745), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n741), .A2(G2067), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT116), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n806), .B(new_n809), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n776), .B(new_n780), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n1001), .A2(G1986), .A3(G290), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT48), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1019), .A2(new_n809), .A3(new_n806), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1002), .B1(new_n1020), .B2(new_n1004), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1002), .A2(new_n876), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1005), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT126), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1002), .A2(new_n780), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT46), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT47), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1018), .A2(new_n1021), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT63), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n506), .A2(new_n999), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n497), .B2(new_n505), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT115), .B1(new_n478), .B2(new_n993), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n1041));
  NOR4_X1   g616(.A1(new_n1041), .A2(new_n467), .A3(new_n995), .A4(new_n992), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1039), .A2(new_n1043), .A3(G2090), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(G1384), .C1(new_n497), .C2(new_n505), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1000), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1971), .B1(new_n1047), .B2(new_n998), .ZN(new_n1048));
  OAI21_X1  g623(.A(G8), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(G166), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n544), .B1(new_n520), .B2(new_n526), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1050), .C1(new_n1054), .C2(new_n518), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n532), .A2(G86), .B1(new_n534), .B2(G48), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n786), .A3(new_n583), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1036), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT121), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(new_n1066), .A3(new_n1069), .A4(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n577), .A2(G1976), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(G8), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT120), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1068), .A2(new_n1070), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1066), .A2(KEYINPUT119), .A3(G8), .A4(new_n1071), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(KEYINPUT52), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1053), .A2(new_n1082), .A3(new_n1055), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(G8), .C1(new_n1044), .C2(new_n1048), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1057), .A2(new_n1077), .A3(new_n1081), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1034), .A2(new_n1045), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1091), .B2(new_n1043), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT50), .B(G1384), .C1(new_n497), .C2(new_n505), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n998), .A3(new_n752), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(G8), .A3(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1033), .B1(new_n1087), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1086), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1056), .ZN(new_n1101));
  INV_X1    g676(.A(G1971), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1091), .B2(new_n1043), .ZN(new_n1103));
  INV_X1    g678(.A(G2090), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1095), .A2(new_n998), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1106), .B2(G8), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1081), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G168), .A2(G8), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1033), .B(new_n1113), .C1(new_n1092), .C2(new_n1096), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1057), .A2(new_n1086), .A3(new_n1114), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1099), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n577), .A2(new_n1074), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT122), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1060), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1052), .B1(new_n998), .B2(new_n1036), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1124), .B1(new_n1111), .B2(new_n1100), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1119), .A2(KEYINPUT124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT124), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1092), .A2(G168), .A3(new_n1096), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(G168), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1132), .A3(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1131), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1047), .A2(new_n998), .A3(new_n727), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1095), .A2(new_n998), .ZN(new_n1140));
  INV_X1    g715(.A(G1961), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1138), .A2(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1139), .A2(G2078), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1047), .A2(new_n998), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(G301), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1087), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1135), .A2(new_n1137), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1047), .A2(new_n998), .A3(new_n780), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT58), .B(G1341), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n1066), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n850), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1348), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n998), .A2(new_n745), .A3(new_n1036), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n852), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1156), .A2(new_n612), .A3(KEYINPUT60), .A4(new_n1157), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n565), .B2(new_n569), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G1956), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT56), .B(G2072), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1047), .A2(new_n998), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1165), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1169), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(KEYINPUT61), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1154), .A2(new_n1164), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n852), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1180), .B1(new_n1183), .B2(new_n1175), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(G301), .A4(new_n1144), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1142), .A2(new_n1190), .A3(G301), .A4(new_n1144), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT54), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1047), .A2(G40), .A3(new_n478), .A4(new_n1143), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1142), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1195), .B2(G171), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1087), .ZN(new_n1198));
  AND4_X1   g773(.A1(G301), .A2(new_n1186), .A3(new_n1187), .A4(new_n1194), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1193), .B1(new_n1145), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1134), .A4(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1148), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1126), .A2(new_n1127), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(G290), .B(new_n811), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1012), .B1(new_n1001), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1032), .B1(new_n1203), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g781(.A1(new_n912), .A2(new_n906), .A3(new_n905), .ZN(new_n1208));
  INV_X1    g782(.A(new_n666), .ZN(new_n1209));
  OR2_X1    g783(.A1(G227), .A2(new_n458), .ZN(new_n1210));
  NOR3_X1   g784(.A1(G229), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n1208), .A2(new_n987), .A3(new_n1211), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


