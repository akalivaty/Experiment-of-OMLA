

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  NOR2_X1 U321 ( .A1(n508), .A2(n487), .ZN(n376) );
  XNOR2_X1 U322 ( .A(n348), .B(n289), .ZN(n349) );
  XNOR2_X1 U323 ( .A(KEYINPUT38), .B(n443), .ZN(n464) );
  INV_X1 U324 ( .A(n546), .ZN(n508) );
  AND2_X1 U325 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U326 ( .A(n344), .B(G127GAT), .Z(n290) );
  INV_X1 U327 ( .A(KEYINPUT96), .ZN(n377) );
  XNOR2_X1 U328 ( .A(n377), .B(KEYINPUT25), .ZN(n378) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U330 ( .A(n402), .B(n349), .ZN(n353) );
  INV_X1 U331 ( .A(G43GAT), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n444), .B(KEYINPUT40), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n446), .B(n445), .ZN(G1330GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n292) );
  NAND2_X1 U335 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U337 ( .A(n293), .B(KEYINPUT73), .Z(n298) );
  XOR2_X1 U338 ( .A(G29GAT), .B(G43GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n424) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n296), .B(G218GAT), .ZN(n369) );
  XNOR2_X1 U343 ( .A(n424), .B(n369), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(G92GAT), .Z(n300) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U348 ( .A(n302), .B(n301), .Z(n304) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G162GAT), .Z(n325) );
  XOR2_X1 U350 ( .A(G99GAT), .B(G85GAT), .Z(n428) );
  XNOR2_X1 U351 ( .A(n325), .B(n428), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n556) );
  XOR2_X1 U353 ( .A(KEYINPUT36), .B(KEYINPUT99), .Z(n305) );
  XNOR2_X1 U354 ( .A(n556), .B(n305), .ZN(n578) );
  XOR2_X1 U355 ( .A(G64GAT), .B(G78GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(G8GAT), .B(G211GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n321) );
  XOR2_X1 U358 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n309) );
  XNOR2_X1 U359 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U361 ( .A(G22GAT), .B(G155GAT), .Z(n324) );
  XOR2_X1 U362 ( .A(n324), .B(G127GAT), .Z(n311) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G1GAT), .Z(n421) );
  XNOR2_X1 U364 ( .A(n421), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U366 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n316), .B(KEYINPUT74), .Z(n319) );
  XNOR2_X1 U370 ( .A(G71GAT), .B(G57GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n317), .B(KEYINPUT13), .ZN(n427) );
  XNOR2_X1 U372 ( .A(n427), .B(KEYINPUT14), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n553) );
  INV_X1 U375 ( .A(n553), .ZN(n574) );
  XOR2_X1 U376 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n323) );
  XNOR2_X1 U377 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT22), .B(G218GAT), .Z(n327) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U383 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n334) );
  XOR2_X1 U385 ( .A(KEYINPUT86), .B(KEYINPUT3), .Z(n333) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n393) );
  XOR2_X1 U388 ( .A(n334), .B(n393), .Z(n341) );
  XOR2_X1 U389 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U392 ( .A(G197GAT), .B(n337), .Z(n370) );
  XOR2_X1 U393 ( .A(G78GAT), .B(G148GAT), .Z(n339) );
  XNOR2_X1 U394 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n438) );
  XNOR2_X1 U396 ( .A(n370), .B(n438), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n542) );
  XOR2_X1 U398 ( .A(KEYINPUT78), .B(KEYINPUT0), .Z(n343) );
  XNOR2_X1 U399 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U401 ( .A(G113GAT), .B(G120GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n290), .B(n345), .ZN(n402) );
  XOR2_X1 U403 ( .A(G190GAT), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(G43GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n351) );
  XNOR2_X1 U407 ( .A(G15GAT), .B(G99GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U409 ( .A(n353), .B(n352), .Z(n361) );
  XOR2_X1 U410 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n355) );
  XNOR2_X1 U411 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(KEYINPUT17), .B(n356), .Z(n371) );
  XOR2_X1 U414 ( .A(G176GAT), .B(KEYINPUT20), .Z(n358) );
  XNOR2_X1 U415 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n371), .B(n359), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n546) );
  XOR2_X1 U419 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XOR2_X1 U420 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n363) );
  XNOR2_X1 U421 ( .A(KEYINPUT95), .B(KEYINPUT93), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U423 ( .A(n423), .B(n364), .Z(n366) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n375) );
  XOR2_X1 U426 ( .A(G64GAT), .B(G92GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(G176GAT), .B(G204GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n437) );
  XOR2_X1 U429 ( .A(n369), .B(n437), .Z(n373) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n536) );
  INV_X1 U433 ( .A(n536), .ZN(n487) );
  NOR2_X1 U434 ( .A1(n542), .A2(n376), .ZN(n379) );
  XOR2_X1 U435 ( .A(n536), .B(KEYINPUT27), .Z(n404) );
  NAND2_X1 U436 ( .A1(n508), .A2(n542), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n380), .B(KEYINPUT26), .ZN(n565) );
  NOR2_X1 U438 ( .A1(n404), .A2(n565), .ZN(n381) );
  NOR2_X1 U439 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n383), .B(KEYINPUT97), .ZN(n403) );
  XOR2_X1 U441 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n385) );
  NAND2_X1 U442 ( .A1(G225GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT5), .B(n386), .ZN(n400) );
  XOR2_X1 U445 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n388) );
  XNOR2_X1 U446 ( .A(G155GAT), .B(KEYINPUT88), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U448 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n390) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(G57GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U451 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U452 ( .A(G85GAT), .B(G162GAT), .Z(n395) );
  XNOR2_X1 U453 ( .A(G29GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(G148GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n540) );
  INV_X1 U459 ( .A(n540), .ZN(n468) );
  AND2_X1 U460 ( .A1(n403), .A2(n540), .ZN(n407) );
  XOR2_X1 U461 ( .A(n542), .B(KEYINPUT28), .Z(n510) );
  NOR2_X1 U462 ( .A1(n404), .A2(n540), .ZN(n507) );
  NAND2_X1 U463 ( .A1(n510), .A2(n507), .ZN(n405) );
  NOR2_X1 U464 ( .A1(n546), .A2(n405), .ZN(n406) );
  NOR2_X1 U465 ( .A1(n407), .A2(n406), .ZN(n449) );
  NOR2_X1 U466 ( .A1(n574), .A2(n449), .ZN(n408) );
  NAND2_X1 U467 ( .A1(n578), .A2(n408), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n409), .B(KEYINPUT37), .ZN(n482) );
  XOR2_X1 U469 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n411) );
  NAND2_X1 U470 ( .A1(G229GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U472 ( .A(n412), .B(KEYINPUT65), .Z(n420) );
  XOR2_X1 U473 ( .A(G197GAT), .B(G113GAT), .Z(n414) );
  XNOR2_X1 U474 ( .A(G36GAT), .B(G50GAT), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U476 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n416) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(G22GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U481 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n547) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U485 ( .A1(G230GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U487 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n432) );
  XNOR2_X1 U488 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n434) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(KEYINPUT68), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n569) );
  NOR2_X1 U497 ( .A1(n547), .A2(n569), .ZN(n450) );
  NAND2_X1 U498 ( .A1(n482), .A2(n450), .ZN(n443) );
  NOR2_X1 U499 ( .A1(n464), .A2(n508), .ZN(n446) );
  NOR2_X1 U500 ( .A1(n556), .A2(n553), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT16), .B(n447), .Z(n448) );
  NOR2_X1 U502 ( .A1(n449), .A2(n448), .ZN(n466) );
  NAND2_X1 U503 ( .A1(n450), .A2(n466), .ZN(n457) );
  NOR2_X1 U504 ( .A1(n540), .A2(n457), .ZN(n451) );
  XOR2_X1 U505 ( .A(G1GAT), .B(n451), .Z(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT34), .B(n452), .ZN(G1324GAT) );
  NOR2_X1 U507 ( .A1(n487), .A2(n457), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT98), .B(n453), .Z(n454) );
  XNOR2_X1 U509 ( .A(G8GAT), .B(n454), .ZN(G1325GAT) );
  NOR2_X1 U510 ( .A1(n508), .A2(n457), .ZN(n456) );
  XNOR2_X1 U511 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(G1326GAT) );
  NOR2_X1 U513 ( .A1(n510), .A2(n457), .ZN(n458) );
  XOR2_X1 U514 ( .A(G22GAT), .B(n458), .Z(G1327GAT) );
  NOR2_X1 U515 ( .A1(n540), .A2(n464), .ZN(n462) );
  XOR2_X1 U516 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n460) );
  XNOR2_X1 U517 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(G1328GAT) );
  NOR2_X1 U520 ( .A1(n464), .A2(n487), .ZN(n463) );
  XOR2_X1 U521 ( .A(G36GAT), .B(n463), .Z(G1329GAT) );
  NOR2_X1 U522 ( .A1(n510), .A2(n464), .ZN(n465) );
  XOR2_X1 U523 ( .A(G50GAT), .B(n465), .Z(G1331GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n470) );
  INV_X1 U525 ( .A(n547), .ZN(n566) );
  XOR2_X1 U526 ( .A(n569), .B(KEYINPUT41), .Z(n526) );
  INV_X1 U527 ( .A(n526), .ZN(n549) );
  NOR2_X1 U528 ( .A1(n566), .A2(n549), .ZN(n483) );
  NAND2_X1 U529 ( .A1(n483), .A2(n466), .ZN(n467) );
  XOR2_X1 U530 ( .A(KEYINPUT102), .B(n467), .Z(n478) );
  NAND2_X1 U531 ( .A1(n468), .A2(n478), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U533 ( .A(G57GAT), .B(n471), .ZN(G1332GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n473) );
  NAND2_X1 U535 ( .A1(n536), .A2(n478), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U537 ( .A(G64GAT), .B(n474), .ZN(G1333GAT) );
  NAND2_X1 U538 ( .A1(n478), .A2(n546), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n475), .B(KEYINPUT106), .ZN(n476) );
  XNOR2_X1 U540 ( .A(G71GAT), .B(n476), .ZN(G1334GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n480) );
  INV_X1 U542 ( .A(n510), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U545 ( .A(G78GAT), .B(n481), .Z(G1335GAT) );
  NAND2_X1 U546 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT108), .ZN(n491) );
  NOR2_X1 U548 ( .A1(n491), .A2(n540), .ZN(n486) );
  XNOR2_X1 U549 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n486), .B(n485), .ZN(G1336GAT) );
  NOR2_X1 U551 ( .A1(n491), .A2(n487), .ZN(n488) );
  XOR2_X1 U552 ( .A(G92GAT), .B(n488), .Z(G1337GAT) );
  NOR2_X1 U553 ( .A1(n491), .A2(n508), .ZN(n489) );
  XOR2_X1 U554 ( .A(KEYINPUT110), .B(n489), .Z(n490) );
  XNOR2_X1 U555 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  NOR2_X1 U556 ( .A1(n510), .A2(n491), .ZN(n492) );
  XOR2_X1 U557 ( .A(KEYINPUT44), .B(n492), .Z(n493) );
  XNOR2_X1 U558 ( .A(G106GAT), .B(n493), .ZN(G1339GAT) );
  NOR2_X1 U559 ( .A1(n547), .A2(n549), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(KEYINPUT46), .ZN(n495) );
  NOR2_X1 U561 ( .A1(n556), .A2(n495), .ZN(n496) );
  NAND2_X1 U562 ( .A1(n496), .A2(n553), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(KEYINPUT47), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n499) );
  NAND2_X1 U565 ( .A1(n574), .A2(n578), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n499), .B(n498), .ZN(n501) );
  INV_X1 U567 ( .A(n569), .ZN(n500) );
  NAND2_X1 U568 ( .A1(n501), .A2(n500), .ZN(n502) );
  NOR2_X1 U569 ( .A1(n566), .A2(n502), .ZN(n503) );
  NOR2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT48), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT111), .ZN(n535) );
  NAND2_X1 U573 ( .A1(n535), .A2(n507), .ZN(n523) );
  NOR2_X1 U574 ( .A1(n508), .A2(n523), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT112), .B(n509), .ZN(n511) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT113), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n566), .A2(n520), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n515) );
  NAND2_X1 U581 ( .A1(n520), .A2(n526), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G120GAT), .B(n516), .ZN(G1341GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n518) );
  NAND2_X1 U585 ( .A1(n520), .A2(n574), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(G127GAT), .B(n519), .ZN(G1342GAT) );
  XOR2_X1 U588 ( .A(G134GAT), .B(KEYINPUT51), .Z(n522) );
  NAND2_X1 U589 ( .A1(n520), .A2(n556), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1343GAT) );
  XNOR2_X1 U591 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n565), .A2(n523), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n532), .A2(n566), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(G1344GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n528) );
  NAND2_X1 U596 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n530) );
  XOR2_X1 U598 ( .A(G148GAT), .B(KEYINPUT117), .Z(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(G1345GAT) );
  NAND2_X1 U600 ( .A1(n532), .A2(n574), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n531), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U602 ( .A1(n532), .A2(n556), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n533), .B(KEYINPUT118), .ZN(n534) );
  XNOR2_X1 U604 ( .A(G162GAT), .B(n534), .ZN(G1347GAT) );
  NAND2_X1 U605 ( .A1(n536), .A2(n535), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n537), .B(KEYINPUT119), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n564) );
  NOR2_X1 U610 ( .A1(n542), .A2(n564), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n547), .A2(n557), .ZN(n548) );
  XOR2_X1 U615 ( .A(G169GAT), .B(n548), .Z(G1348GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n557), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(n552), .ZN(G1349GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n557), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G183GAT), .B(n555), .ZN(G1350GAT) );
  INV_X1 U623 ( .A(n556), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U625 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(n561), .ZN(G1351GAT) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT124), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(n563), .Z(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U635 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT127), .Z(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

