

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U323 ( .A1(n538), .A2(n460), .ZN(n564) );
  XOR2_X1 U324 ( .A(KEYINPUT40), .B(n507), .Z(n291) );
  INV_X1 U325 ( .A(KEYINPUT31), .ZN(n371) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n414) );
  XNOR2_X1 U327 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U328 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n415), .B(n414), .ZN(n535) );
  XNOR2_X1 U330 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U331 ( .A(n374), .B(n373), .ZN(n378) );
  XNOR2_X1 U332 ( .A(n496), .B(KEYINPUT103), .ZN(n497) );
  NOR2_X1 U333 ( .A1(n477), .A2(n476), .ZN(n494) );
  XNOR2_X1 U334 ( .A(n498), .B(n497), .ZN(n521) );
  XOR2_X1 U335 ( .A(KEYINPUT41), .B(n577), .Z(n554) );
  XOR2_X1 U336 ( .A(n366), .B(n365), .Z(n574) );
  XOR2_X1 U337 ( .A(n470), .B(KEYINPUT28), .Z(n540) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n464) );
  XNOR2_X1 U339 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(G176GAT), .B(KEYINPUT84), .Z(n293) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G113GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U343 ( .A(KEYINPUT83), .B(G99GAT), .Z(n295) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U346 ( .A(KEYINPUT81), .B(KEYINPUT87), .Z(n297) );
  XNOR2_X1 U347 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U350 ( .A(G120GAT), .B(G71GAT), .Z(n370) );
  XOR2_X1 U351 ( .A(G134GAT), .B(KEYINPUT0), .Z(n442) );
  XOR2_X1 U352 ( .A(G15GAT), .B(G127GAT), .Z(n338) );
  XOR2_X1 U353 ( .A(n442), .B(n338), .Z(n301) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n370), .B(n302), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n311) );
  XOR2_X1 U359 ( .A(G183GAT), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U360 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n309) );
  XOR2_X1 U363 ( .A(n310), .B(n309), .Z(n329) );
  XNOR2_X1 U364 ( .A(n311), .B(n329), .ZN(n486) );
  INV_X1 U365 ( .A(n486), .ZN(n538) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G92GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n312), .B(G64GAT), .ZN(n381) );
  XOR2_X1 U368 ( .A(G36GAT), .B(G190GAT), .Z(n388) );
  XNOR2_X1 U369 ( .A(n381), .B(n388), .ZN(n313) );
  AND2_X1 U370 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  NAND2_X1 U371 ( .A1(n313), .A2(n314), .ZN(n318) );
  INV_X1 U372 ( .A(n313), .ZN(n316) );
  INV_X1 U373 ( .A(n314), .ZN(n315) );
  NAND2_X1 U374 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND2_X1 U375 ( .A1(n318), .A2(n317), .ZN(n324) );
  XOR2_X1 U376 ( .A(G204GAT), .B(G211GAT), .Z(n320) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n419) );
  XNOR2_X1 U379 ( .A(n419), .B(KEYINPUT97), .ZN(n322) );
  INV_X1 U380 ( .A(KEYINPUT96), .ZN(n321) );
  XOR2_X1 U381 ( .A(n325), .B(KEYINPUT75), .Z(n327) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G8GAT), .Z(n362) );
  XNOR2_X1 U383 ( .A(n362), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n504) );
  XOR2_X1 U386 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n331) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U389 ( .A(KEYINPUT75), .B(G78GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n351) );
  XOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n337) );
  XNOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT80), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XOR2_X1 U397 ( .A(n427), .B(n338), .Z(n340) );
  XNOR2_X1 U398 ( .A(G183GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n344) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n345), .B(KEYINPUT14), .Z(n349) );
  XOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT66), .Z(n347) );
  XNOR2_X1 U405 ( .A(G57GAT), .B(KEYINPUT67), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n367) );
  XNOR2_X1 U407 ( .A(n367), .B(KEYINPUT76), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n580) );
  XOR2_X1 U410 ( .A(G197GAT), .B(G15GAT), .Z(n353) );
  XNOR2_X1 U411 ( .A(G36GAT), .B(G50GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n366) );
  XOR2_X1 U413 ( .A(G29GAT), .B(G43GAT), .Z(n355) );
  XNOR2_X1 U414 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n401) );
  XOR2_X1 U416 ( .A(n401), .B(KEYINPUT30), .Z(n357) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U419 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n359) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n361), .B(n360), .Z(n364) );
  XOR2_X1 U423 ( .A(G113GAT), .B(G1GAT), .Z(n449) );
  XNOR2_X1 U424 ( .A(n449), .B(n362), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U426 ( .A(G99GAT), .B(G85GAT), .Z(n387) );
  XNOR2_X1 U427 ( .A(n367), .B(n387), .ZN(n369) );
  AND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n370), .B(G204GAT), .ZN(n372) );
  XOR2_X1 U431 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n376) );
  XNOR2_X1 U432 ( .A(KEYINPUT32), .B(KEYINPUT68), .ZN(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G148GAT), .Z(n380) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n423) );
  XNOR2_X1 U438 ( .A(n423), .B(n381), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n577) );
  NAND2_X1 U440 ( .A1(n574), .A2(n554), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT46), .ZN(n404) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n386) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT9), .B(n387), .Z(n390) );
  XNOR2_X1 U446 ( .A(n388), .B(G92GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U451 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n396) );
  XNOR2_X1 U452 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U454 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U455 ( .A(G162GAT), .B(KEYINPUT71), .Z(n400) );
  XNOR2_X1 U456 ( .A(G50GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n420) );
  XNOR2_X1 U458 ( .A(n401), .B(n420), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n478) );
  NAND2_X1 U460 ( .A1(n404), .A2(n478), .ZN(n405) );
  NOR2_X1 U461 ( .A1(n580), .A2(n405), .ZN(n406) );
  XOR2_X1 U462 ( .A(n406), .B(KEYINPUT47), .Z(n413) );
  INV_X1 U463 ( .A(n478), .ZN(n561) );
  XNOR2_X1 U464 ( .A(KEYINPUT36), .B(n561), .ZN(n583) );
  NAND2_X1 U465 ( .A1(n583), .A2(n580), .ZN(n408) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  INV_X1 U468 ( .A(n574), .ZN(n512) );
  NAND2_X1 U469 ( .A1(n409), .A2(n512), .ZN(n410) );
  NOR2_X1 U470 ( .A1(n577), .A2(n410), .ZN(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT114), .B(n411), .ZN(n412) );
  NOR2_X1 U472 ( .A1(n413), .A2(n412), .ZN(n415) );
  NAND2_X1 U473 ( .A1(n504), .A2(n535), .ZN(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n416), .B(KEYINPUT54), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n571) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n433) );
  XOR2_X1 U478 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n422) );
  XNOR2_X1 U479 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n443) );
  XNOR2_X1 U481 ( .A(n423), .B(n443), .ZN(n431) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n470) );
  XOR2_X1 U490 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n435) );
  XNOR2_X1 U491 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n457) );
  XOR2_X1 U493 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n437) );
  XNOR2_X1 U494 ( .A(G148GAT), .B(KEYINPUT91), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U496 ( .A(G57GAT), .B(KEYINPUT92), .Z(n439) );
  XNOR2_X1 U497 ( .A(KEYINPUT95), .B(KEYINPUT6), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n455) );
  XOR2_X1 U500 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U501 ( .A1(G225GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n453) );
  XOR2_X1 U503 ( .A(G162GAT), .B(G155GAT), .Z(n447) );
  XNOR2_X1 U504 ( .A(G120GAT), .B(G127GAT), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U506 ( .A(n448), .B(G85GAT), .Z(n451) );
  XNOR2_X1 U507 ( .A(n449), .B(G29GAT), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n570) );
  INV_X1 U512 ( .A(n570), .ZN(n482) );
  NOR2_X1 U513 ( .A1(n470), .A2(n482), .ZN(n458) );
  AND2_X1 U514 ( .A1(n571), .A2(n458), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT55), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n564), .A2(n554), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NAND2_X1 U520 ( .A1(n561), .A2(n564), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT27), .B(n504), .Z(n472) );
  NOR2_X1 U522 ( .A1(n570), .A2(n472), .ZN(n536) );
  NAND2_X1 U523 ( .A1(n536), .A2(n540), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n486), .A2(n466), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT98), .ZN(n477) );
  AND2_X1 U526 ( .A1(n504), .A2(n486), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n470), .A2(n468), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n469), .Z(n474) );
  NAND2_X1 U529 ( .A1(n538), .A2(n470), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT26), .ZN(n573) );
  NOR2_X1 U531 ( .A1(n573), .A2(n472), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n482), .A2(n475), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n478), .A2(n580), .ZN(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT16), .B(n479), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n494), .A2(n480), .ZN(n513) );
  NOR2_X1 U537 ( .A1(n577), .A2(n512), .ZN(n499) );
  NAND2_X1 U538 ( .A1(n513), .A2(n499), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT99), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n491), .A2(n482), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n504), .A2(n491), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U546 ( .A1(n491), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT101), .Z(n493) );
  INV_X1 U550 ( .A(n540), .ZN(n490) );
  NAND2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  NOR2_X1 U553 ( .A1(n580), .A2(n494), .ZN(n495) );
  NAND2_X1 U554 ( .A1(n583), .A2(n495), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT37), .B(KEYINPUT102), .Z(n496) );
  NAND2_X1 U556 ( .A1(n521), .A2(n499), .ZN(n500) );
  XNOR2_X1 U557 ( .A(n500), .B(KEYINPUT38), .ZN(n501) );
  XNOR2_X1 U558 ( .A(KEYINPUT104), .B(n501), .ZN(n508) );
  NOR2_X1 U559 ( .A1(n570), .A2(n508), .ZN(n502) );
  XNOR2_X1 U560 ( .A(n502), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  INV_X1 U562 ( .A(n504), .ZN(n526) );
  NOR2_X1 U563 ( .A1(n526), .A2(n508), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(G1329GAT) );
  NOR2_X1 U566 ( .A1(n538), .A2(n508), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n291), .ZN(G1330GAT) );
  NOR2_X1 U568 ( .A1(n540), .A2(n508), .ZN(n509) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n511) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n515) );
  AND2_X1 U573 ( .A1(n512), .A2(n554), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n513), .A2(n522), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n570), .A2(n518), .ZN(n514) );
  XOR2_X1 U576 ( .A(n515), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n526), .A2(n518), .ZN(n516) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n538), .A2(n518), .ZN(n517) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n540), .A2(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n570), .A2(n532), .ZN(n524) );
  XNOR2_X1 U586 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n527), .Z(n528) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n538), .A2(n532), .ZN(n529) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n534) );
  NOR2_X1 U597 ( .A1(n540), .A2(n532), .ZN(n533) );
  XOR2_X1 U598 ( .A(n534), .B(n533), .Z(G1339GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT116), .ZN(n551) );
  NOR2_X1 U601 ( .A1(n551), .A2(n538), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U603 ( .A(KEYINPUT117), .B(n541), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n548), .A2(n574), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n544) );
  NAND2_X1 U607 ( .A1(n548), .A2(n554), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n548), .A2(n580), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U614 ( .A1(n548), .A2(n561), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT119), .Z(n553) );
  NOR2_X1 U617 ( .A1(n551), .A2(n573), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n574), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U622 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n580), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n574), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .Z(n566) );
  NAND2_X1 U632 ( .A1(n564), .A2(n580), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(n569), .Z(n576) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

