//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT81), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G78gat), .B(G106gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT22), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G211gat), .A2(G218gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n210), .B(new_n211), .C1(new_n209), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(KEYINPUT22), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n209), .A2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n216), .B2(KEYINPUT71), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(KEYINPUT71), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT77), .B(G141gat), .Z(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G141gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n221), .A2(new_n224), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT74), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n232), .A2(new_n233), .B1(G155gat), .B2(G162gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n235));
  XOR2_X1   g034(.A(G141gat), .B(G148gat), .Z(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT75), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT75), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n222), .A2(G148gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n224), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n234), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT76), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n243), .B(new_n234), .C1(new_n237), .C2(new_n240), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n230), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n219), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n213), .A2(new_n216), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n248), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n245), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n206), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT80), .B(new_n206), .C1(new_n249), .C2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT3), .B1(new_n219), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(G228gat), .B(G233gat), .C1(new_n259), .C2(new_n245), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(new_n249), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G22gat), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n205), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n257), .B2(new_n262), .ZN(new_n268));
  AOI211_X1 g067(.A(G22gat), .B(new_n261), .C1(new_n255), .C2(new_n256), .ZN(new_n269));
  INV_X1    g068(.A(new_n205), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n204), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n266), .A3(new_n205), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n203), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  INV_X1    g076(.A(G226gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT65), .Z(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n281), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n283), .B(KEYINPUT66), .Z(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n287), .C1(KEYINPUT26), .C2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n292), .B2(KEYINPUT67), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  MUX2_X1   g097(.A(KEYINPUT24), .B(new_n298), .S(new_n295), .Z(new_n299));
  AND2_X1   g098(.A1(new_n299), .A2(new_n281), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(new_n283), .B2(KEYINPUT23), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(new_n283), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n283), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n303), .B2(new_n302), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n300), .B(new_n309), .C1(new_n302), .C2(new_n288), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n289), .A2(new_n297), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI221_X1 g110(.A(new_n277), .B1(new_n278), .B2(new_n279), .C1(new_n311), .C2(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n297), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n310), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n278), .A2(new_n279), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n316), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n312), .A2(new_n317), .A3(new_n319), .A4(new_n219), .ZN(new_n320));
  INV_X1    g119(.A(new_n248), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  INV_X1    g122(.A(new_n219), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G64gat), .B(G92gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n320), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(KEYINPUT30), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n330), .A2(KEYINPUT30), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(new_n325), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n328), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(G127gat), .B2(G134gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(G127gat), .B2(G134gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT1), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n338), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n247), .B(new_n342), .C1(new_n343), .C2(new_n245), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n245), .A2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(new_n345), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n351));
  INV_X1    g150(.A(new_n245), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n342), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(new_n345), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(KEYINPUT5), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT79), .A3(new_n350), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  INV_X1    g165(.A(new_n364), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n357), .A2(new_n367), .A3(new_n359), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n367), .A4(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n335), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n311), .B(new_n342), .ZN(new_n372));
  AND2_X1   g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT34), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n377), .A3(new_n378), .A4(new_n374), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT70), .B1(new_n375), .B2(KEYINPUT34), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  XOR2_X1   g181(.A(G15gat), .B(G43gat), .Z(new_n383));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI221_X1 g185(.A(KEYINPUT32), .B1(new_n382), .B2(new_n386), .C1(new_n372), .C2(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n382), .B1(new_n372), .B2(new_n374), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT32), .B1(new_n372), .B2(new_n374), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(new_n381), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n387), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n381), .A2(new_n379), .A3(new_n376), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n276), .A2(new_n371), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT35), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n370), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n370), .A2(new_n399), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n369), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n335), .A2(KEYINPUT35), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n272), .B2(new_n275), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT36), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT36), .B1(new_n391), .B2(new_n394), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n275), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n203), .B1(new_n273), .B2(new_n274), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n369), .A2(new_n370), .ZN(new_n413));
  INV_X1    g212(.A(new_n335), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n348), .A2(new_n349), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n345), .B1(new_n417), .B2(new_n344), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT39), .B1(new_n354), .B2(new_n355), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT39), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n364), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT40), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(new_n335), .A3(new_n368), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT38), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT37), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n320), .A2(new_n325), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n430), .A2(new_n328), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n333), .A2(KEYINPUT37), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n323), .B2(new_n219), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n312), .A2(new_n317), .A3(new_n319), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(new_n219), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(new_n430), .A3(new_n428), .A4(new_n328), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n330), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n276), .B(new_n427), .C1(new_n402), .C2(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n398), .A2(new_n406), .B1(new_n416), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G1gat), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n265), .A2(G15gat), .ZN(new_n444));
  INV_X1    g243(.A(G15gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G22gat), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n447), .A2(G8gat), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G8gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G1gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT86), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(G8gat), .B1(new_n447), .B2(new_n448), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n453), .A3(new_n450), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g260(.A(G43gat), .ZN(new_n462));
  INV_X1    g261(.A(G50gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G43gat), .A2(G50gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT15), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT84), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(G29gat), .A3(G36gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT14), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT14), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(G29gat), .B2(G36gat), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n461), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n481), .A2(KEYINPUT85), .A3(new_n467), .A4(new_n469), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(KEYINPUT15), .A3(new_n466), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n460), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n449), .A2(new_n454), .A3(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n458), .B1(new_n456), .B2(new_n457), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n484), .B(new_n490), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT13), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n491), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n490), .B1(new_n460), .B2(new_n484), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n497), .A2(new_n498), .B1(new_n484), .B2(new_n460), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n494), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n489), .A2(new_n491), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n480), .A2(new_n482), .A3(new_n505), .A4(new_n483), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n456), .A2(new_n457), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(new_n493), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n496), .A2(new_n501), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n503), .A2(new_n509), .A3(KEYINPUT18), .A4(new_n493), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT88), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n489), .A2(new_n491), .B1(new_n507), .B2(new_n508), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT18), .A4(new_n493), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G169gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G197gat), .ZN(new_n522));
  INV_X1    g321(.A(G169gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n520), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G197gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT12), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n511), .A2(new_n517), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n528), .B2(new_n530), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n511), .B2(new_n517), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n441), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G183gat), .B(G211gat), .Z(new_n540));
  XOR2_X1   g339(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G57gat), .B(G64gat), .Z(new_n543));
  OR2_X1    g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n543), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n545), .B(new_n544), .C1(new_n552), .C2(new_n548), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT21), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n542), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n460), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n551), .A2(KEYINPUT21), .A3(new_n553), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n559), .A3(new_n542), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n561), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n540), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n565), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n562), .B(new_n563), .C1(new_n569), .C2(new_n560), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n571));
  INV_X1    g370(.A(new_n540), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT91), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G92gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G99gat), .ZN(new_n582));
  INV_X1    g381(.A(G106gat), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT8), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(KEYINPUT92), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n575), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n581), .A2(KEYINPUT92), .A3(new_n584), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT92), .B1(new_n581), .B2(new_n584), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n575), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n484), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n504), .B2(new_n506), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n601), .B2(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n606), .A2(new_n607), .A3(new_n614), .A4(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n574), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n574), .A2(KEYINPUT94), .A3(new_n618), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n551), .A2(new_n624), .A3(new_n553), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n592), .B2(new_n596), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n628));
  INV_X1    g427(.A(new_n575), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n551), .A2(new_n553), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT95), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n630), .A2(new_n595), .A3(new_n632), .A4(new_n625), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n595), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT96), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n630), .A2(new_n636), .A3(new_n639), .A4(new_n595), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n634), .A2(new_n635), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n623), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n638), .A2(new_n640), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT10), .B1(new_n627), .B2(new_n633), .ZN(new_n646));
  OAI211_X1 g445(.A(KEYINPUT97), .B(new_n642), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n627), .A2(new_n643), .A3(new_n633), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n644), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT98), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n644), .A2(new_n647), .A3(new_n656), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n646), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n640), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n643), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n652), .B1(new_n661), .B2(new_n649), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n621), .A2(new_n622), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n539), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n413), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n442), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n414), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(G8gat), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(KEYINPUT101), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n671), .B2(new_n672), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n678));
  OAI211_X1 g477(.A(new_n673), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(new_n409), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n667), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n396), .A2(new_n445), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n667), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n276), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR3_X1   g485(.A1(new_n574), .A2(new_n663), .A3(new_n618), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n539), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(G29gat), .A3(new_n413), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n441), .B2(new_n618), .ZN(new_n692));
  INV_X1    g491(.A(new_n618), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n416), .A2(new_n440), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n397), .A2(KEYINPUT35), .B1(new_n405), .B2(new_n404), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT44), .B(new_n693), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n574), .B(KEYINPUT103), .ZN(new_n698));
  INV_X1    g497(.A(new_n537), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n511), .A2(new_n517), .A3(new_n531), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT102), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n532), .A2(new_n537), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n698), .A2(new_n664), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n413), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n707), .ZN(G1328gat));
  NOR3_X1   g507(.A1(new_n688), .A2(G36gat), .A3(new_n414), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n706), .B2(new_n414), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(new_n462), .B1(new_n688), .B2(new_n395), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n409), .A2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g515(.A(new_n463), .B1(new_n688), .B2(new_n276), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n412), .A2(G50gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n706), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g519(.A1(new_n621), .A2(new_n622), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n441), .A2(new_n721), .A3(new_n664), .A4(new_n704), .ZN(new_n722));
  INV_X1    g521(.A(new_n413), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT104), .B(G57gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n335), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n728), .B2(new_n727), .ZN(G1333gat));
  NAND3_X1  g530(.A1(new_n722), .A2(G71gat), .A3(new_n409), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n722), .A2(new_n396), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n734), .B(new_n735), .C1(G71gat), .C2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n412), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n704), .A2(new_n574), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n663), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT107), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n697), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n413), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n693), .B(new_n742), .C1(new_n694), .C2(new_n695), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n398), .A2(new_n406), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n416), .A2(new_n440), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n742), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n664), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n580), .A3(new_n723), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n746), .A2(new_n755), .ZN(G1336gat));
  NAND2_X1  g555(.A1(new_n335), .A2(new_n576), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n692), .A2(new_n696), .A3(new_n335), .A4(new_n744), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n577), .A2(new_n579), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(KEYINPUT108), .A3(new_n762), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n759), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT52), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(KEYINPUT52), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n764), .B1(new_n770), .B2(new_n771), .ZN(G1337gat));
  NOR3_X1   g571(.A1(new_n745), .A2(new_n582), .A3(new_n680), .ZN(new_n773));
  AOI21_X1  g572(.A(G99gat), .B1(new_n754), .B2(new_n396), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1338gat));
  OAI21_X1  g574(.A(G106gat), .B1(new_n745), .B2(new_n276), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n749), .A2(new_n753), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(new_n583), .A3(new_n412), .A4(new_n663), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n665), .A2(new_n704), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n499), .A2(new_n494), .B1(new_n514), .B2(new_n493), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n527), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n700), .A2(new_n616), .A3(new_n617), .A4(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n641), .B2(new_n643), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n644), .A2(new_n786), .A3(new_n647), .ZN(new_n787));
  INV_X1    g586(.A(new_n652), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n661), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n658), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n658), .B2(new_n795), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n784), .B(new_n793), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n700), .A2(new_n783), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n663), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n793), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n658), .A2(new_n795), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT111), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(new_n796), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n802), .B1(new_n806), .B2(new_n704), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n799), .B1(new_n807), .B2(new_n693), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n781), .B1(new_n808), .B2(new_n698), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n413), .A2(new_n335), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR4_X1   g610(.A1(new_n809), .A2(new_n395), .A3(new_n412), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n704), .ZN(new_n813));
  INV_X1    g612(.A(new_n538), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(G113gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(G1340gat));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n663), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(G120gat), .ZN(G1341gat));
  INV_X1    g617(.A(new_n812), .ZN(new_n819));
  INV_X1    g618(.A(G127gat), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n698), .ZN(new_n821));
  INV_X1    g620(.A(new_n574), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(G127gat), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT112), .B1(new_n819), .B2(new_n822), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n693), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n828), .A2(KEYINPUT113), .A3(G134gat), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(new_n828), .B2(G134gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n831), .B2(KEYINPUT56), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n833), .A4(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n831), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n828), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n811), .A2(new_n409), .ZN(new_n838));
  INV_X1    g637(.A(new_n809), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n839), .B2(new_n412), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n412), .A2(KEYINPUT57), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT115), .B1(new_n791), .B2(new_n792), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(KEYINPUT55), .C1(new_n787), .C2(new_n790), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n658), .B(new_n795), .C1(new_n532), .C2(new_n537), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n801), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n801), .B(new_n849), .C1(new_n845), .C2(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n618), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n799), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n822), .ZN(new_n853));
  INV_X1    g652(.A(new_n781), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n841), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n838), .B1(new_n840), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n220), .B1(new_n857), .B2(new_n704), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n809), .A2(new_n811), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n409), .A2(new_n276), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n538), .A2(G141gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n220), .B1(new_n857), .B2(new_n814), .ZN(new_n866));
  INV_X1    g665(.A(new_n863), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n864), .A2(new_n865), .B1(new_n866), .B2(new_n868), .ZN(G1344gat));
  NOR4_X1   g668(.A1(new_n413), .A2(G148gat), .A3(new_n335), .A4(new_n664), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n839), .A2(new_n860), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n666), .A2(new_n538), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n853), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n799), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n693), .B1(new_n847), .B2(KEYINPUT116), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n850), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n873), .B(new_n874), .C1(new_n878), .C2(new_n574), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n276), .A2(KEYINPUT57), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n809), .B2(new_n276), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n663), .A3(new_n838), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n872), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(G148gat), .C1(new_n856), .C2(new_n664), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n885), .B2(KEYINPUT119), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n871), .B1(new_n886), .B2(new_n889), .ZN(G1345gat));
  NOR3_X1   g689(.A1(new_n856), .A2(new_n226), .A3(new_n698), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n861), .A2(KEYINPUT120), .A3(new_n822), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(G155gat), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT120), .B1(new_n861), .B2(new_n822), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n856), .B2(new_n618), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n862), .A2(new_n227), .A3(new_n693), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n809), .A2(new_n723), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n405), .A2(new_n335), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n523), .A3(new_n538), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT121), .B1(new_n809), .B2(new_n723), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n704), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(new_n523), .ZN(G1348gat));
  INV_X1    g709(.A(G176gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n911), .A3(new_n663), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n902), .B2(new_n664), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n290), .A3(new_n574), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n902), .B2(new_n698), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n908), .A2(new_n291), .A3(new_n693), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  INV_X1    g720(.A(new_n902), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n693), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(G190gat), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT61), .B(new_n291), .C1(new_n922), .C2(new_n693), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  AND4_X1   g725(.A1(new_n335), .A2(new_n905), .A3(new_n860), .A4(new_n906), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n704), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n409), .A2(new_n723), .A3(new_n414), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n883), .B1(new_n875), .B2(new_n881), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(KEYINPUT123), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(new_n883), .C1(new_n875), .C2(new_n881), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n538), .A2(new_n525), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  XNOR2_X1  g736(.A(KEYINPUT124), .B(G204gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n664), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n927), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT62), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n935), .A2(new_n663), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n207), .A3(new_n574), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n882), .A2(new_n574), .A3(new_n883), .A4(new_n929), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n693), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n208), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n952), .A2(KEYINPUT125), .A3(new_n934), .A4(new_n929), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n618), .A2(new_n208), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT125), .B1(new_n932), .B2(new_n934), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n951), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


