//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G155gat), .B(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G134gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G127gat), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G120gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n230), .B2(new_n232), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n228), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n230), .ZN(new_n243));
  INV_X1    g042(.A(new_n228), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n245), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n250));
  NAND3_X1  g049(.A1(new_n213), .A2(new_n222), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n213), .A2(new_n222), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n223), .A2(new_n238), .A3(KEYINPUT4), .A4(new_n245), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n248), .A2(new_n254), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n252), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n246), .ZN(new_n261));
  INV_X1    g060(.A(new_n255), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G120gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT1), .B1(new_n265), .B2(new_n233), .ZN(new_n266));
  INV_X1    g065(.A(new_n237), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n244), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n225), .A2(new_n227), .A3(new_n235), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n230), .B2(new_n242), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n268), .A2(new_n252), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n238), .A2(new_n245), .B1(new_n213), .B2(new_n222), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(KEYINPUT75), .B2(new_n257), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n206), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n263), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n205), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT76), .B1(new_n282), .B2(KEYINPUT6), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n205), .A3(new_n281), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT6), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G211gat), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G218gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G211gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n304), .B2(KEYINPUT22), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT69), .B(G211gat), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT70), .B(new_n306), .C1(new_n307), .C2(new_n293), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G197gat), .ZN(new_n310));
  INV_X1    g109(.A(G204gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n299), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  AOI211_X1 g118(.A(new_n298), .B(new_n317), .C1(new_n305), .C2(new_n308), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT24), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT25), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n326), .A2(new_n332), .A3(new_n337), .A4(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G183gat), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT64), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT64), .B1(new_n345), .B2(new_n347), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n334), .A2(KEYINPUT28), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT65), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT65), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n336), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n342), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n323), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n356), .A2(new_n358), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n324), .B1(new_n364), .B2(new_n355), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n347), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT64), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n351), .ZN(new_n370));
  INV_X1    g169(.A(new_n344), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n365), .A2(new_n372), .B1(new_n340), .B2(new_n341), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(new_n322), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT72), .B1(new_n363), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT72), .B1(new_n361), .B2(new_n323), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n321), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT73), .B1(new_n373), .B2(new_n322), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n380), .A3(new_n323), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n322), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n382), .A2(new_n321), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n292), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n321), .A3(new_n383), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n361), .A2(new_n323), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n376), .B1(new_n388), .B2(KEYINPUT72), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n386), .B(new_n291), .C1(new_n389), .C2(new_n321), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(KEYINPUT30), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n378), .A2(new_n384), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n291), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n288), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n288), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(G22gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n309), .A2(new_n318), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n298), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n309), .A2(new_n299), .A3(new_n318), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n362), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n223), .B1(new_n406), .B2(new_n250), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n321), .B1(new_n362), .B2(new_n251), .ZN(new_n408));
  INV_X1    g207(.A(G228gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT3), .B1(new_n406), .B2(KEYINPUT78), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT29), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n223), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n421), .B2(KEYINPUT79), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n406), .A2(KEYINPUT78), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT79), .B(new_n252), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n411), .B(new_n415), .C1(new_n422), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n252), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n426), .A3(new_n416), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n415), .B1(new_n433), .B2(new_n411), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n402), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n411), .B1(new_n422), .B2(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n414), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n401), .A3(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n400), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n276), .A2(new_n278), .A3(new_n284), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(new_n287), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n291), .B1(new_n392), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT37), .B1(new_n378), .B2(new_n384), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n389), .A2(new_n321), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n363), .B1(new_n379), .B2(new_n381), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT83), .B1(new_n450), .B2(new_n321), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n321), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT37), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n446), .B1(new_n454), .B2(new_n445), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n390), .B(new_n443), .C1(new_n448), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n248), .A2(new_n254), .A3(new_n256), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT81), .B(KEYINPUT39), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n262), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n206), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT82), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n262), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(KEYINPUT39), .C1(new_n262), .C2(new_n261), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n286), .B1(new_n464), .B2(KEYINPUT40), .ZN(new_n465));
  INV_X1    g264(.A(new_n395), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n466), .C1(KEYINPUT40), .C2(new_n464), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n456), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n361), .A2(new_n238), .A3(new_n245), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n373), .A2(new_n249), .ZN(new_n470));
  INV_X1    g269(.A(G227gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n410), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G43gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n473), .B(KEYINPUT32), .C1(new_n480), .C2(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n469), .A2(new_n470), .ZN(new_n484));
  INV_X1    g283(.A(new_n472), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(KEYINPUT34), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(KEYINPUT34), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n482), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n482), .B2(new_n483), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n440), .A2(new_n468), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n435), .A2(new_n438), .A3(new_n492), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT35), .B1(new_n400), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n466), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n498), .A2(KEYINPUT85), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(KEYINPUT35), .C1(new_n400), .C2(new_n497), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n507), .A2(KEYINPUT89), .B1(G43gat), .B2(G50gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(KEYINPUT89), .B2(new_n507), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT90), .B(G50gat), .Z(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT88), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n506), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(G8gat), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n529), .ZN(new_n534));
  INV_X1    g333(.A(new_n521), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT87), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G113gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n214), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n529), .B(new_n521), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n537), .B(KEYINPUT13), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n538), .B2(new_n539), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT93), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n551), .C1(new_n538), .C2(new_n539), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n540), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n547), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT94), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n553), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n504), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT98), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n524), .A2(new_n532), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  AND2_X1   g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n580), .A2(new_n535), .B1(KEYINPUT41), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n585), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n593), .B2(new_n592), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT96), .ZN(new_n601));
  INV_X1    g400(.A(new_n591), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n599), .B2(KEYINPUT96), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(new_n596), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n226), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n534), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n575), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n569), .A2(KEYINPUT99), .A3(new_n570), .A4(new_n574), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n566), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT100), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n606), .A3(new_n576), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n578), .A2(new_n605), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT101), .ZN(new_n629));
  XOR2_X1   g428(.A(G120gat), .B(G148gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT102), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT103), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n624), .A2(new_n635), .A3(new_n625), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n578), .A2(new_n635), .A3(new_n605), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n627), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n629), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n634), .B1(new_n629), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n618), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n564), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n288), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n466), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT104), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT42), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(G8gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT105), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n644), .B2(new_n495), .ZN(new_n656));
  INV_X1    g455(.A(new_n492), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n644), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n441), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n617), .ZN(new_n663));
  INV_X1    g462(.A(new_n642), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n590), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n564), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G29gat), .A3(new_n288), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n504), .B2(new_n590), .ZN(new_n672));
  AOI221_X4 g471(.A(KEYINPUT77), .B1(new_n391), .B2(new_n394), .C1(new_n285), .C2(new_n287), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n398), .B1(new_n288), .B2(new_n395), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n497), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT35), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT85), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n499), .A2(new_n500), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n503), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n440), .A2(new_n468), .A3(new_n495), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n590), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n672), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n665), .A2(new_n563), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n288), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n686), .ZN(G1328gat));
  NOR3_X1   g486(.A1(new_n667), .A2(G36gat), .A3(new_n395), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT46), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n685), .B2(new_n395), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1329gat));
  OAI21_X1  g490(.A(new_n510), .B1(new_n667), .B2(new_n657), .ZN(new_n692));
  INV_X1    g491(.A(new_n495), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g495(.A1(new_n564), .A2(new_n439), .A3(new_n666), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n697), .A2(new_n511), .B1(new_n698), .B2(KEYINPUT48), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n441), .A2(new_n511), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n685), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(KEYINPUT48), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n701), .B(new_n702), .Z(G1331gat));
  INV_X1    g502(.A(new_n553), .ZN(new_n704));
  INV_X1    g503(.A(new_n562), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n561), .B1(new_n557), .B2(new_n558), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OR4_X1    g506(.A1(new_n504), .A2(new_n707), .A3(new_n618), .A4(new_n664), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n288), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n599), .ZN(G1332gat));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n395), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n708), .B2(new_n495), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n657), .A2(G71gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n708), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1334gat));
  NOR2_X1   g519(.A1(new_n708), .A2(new_n441), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT109), .B(G78gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n617), .A3(new_n664), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n683), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n288), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n617), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n681), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT51), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n681), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n642), .A2(new_n572), .A3(new_n646), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n726), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT110), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n725), .B2(new_n395), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n664), .A2(G92gat), .A3(new_n395), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n679), .A2(new_n680), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n730), .A2(KEYINPUT111), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n742), .A2(new_n589), .A3(new_n727), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n681), .B2(new_n727), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n747), .B2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n725), .B2(new_n495), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n664), .A2(G99gat), .A3(new_n657), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n733), .B2(new_n751), .ZN(G1338gat));
  NOR3_X1   g551(.A1(new_n664), .A2(G106gat), .A3(new_n441), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n744), .B2(new_n745), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n672), .A2(new_n682), .A3(new_n439), .A4(new_n724), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n758), .A3(G106gat), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT114), .B(new_n753), .C1(new_n744), .C2(new_n745), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n757), .B2(G106gat), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT53), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n732), .A2(new_n753), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n757), .A2(G106gat), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n763), .A2(new_n767), .A3(KEYINPUT116), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1339gat));
  INV_X1    g571(.A(new_n639), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n636), .A2(new_n627), .A3(new_n638), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n634), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n639), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n640), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n533), .A2(new_n536), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n785), .A2(new_n537), .B1(new_n549), .B2(new_n550), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n553), .B1(new_n546), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n589), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n707), .A2(new_n784), .B1(new_n642), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n589), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n790), .A2(new_n663), .B1(new_n563), .B2(new_n643), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n439), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n646), .A2(new_n395), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n657), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n563), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n791), .A2(new_n288), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n499), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n707), .A2(new_n239), .A3(new_n241), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT117), .Z(G1340gat));
  NOR3_X1   g600(.A1(new_n795), .A2(new_n229), .A3(new_n664), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n499), .A3(new_n642), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n229), .B2(new_n803), .ZN(G1341gat));
  OAI21_X1  g603(.A(G127gat), .B1(new_n795), .B2(new_n663), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n617), .A2(new_n226), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n798), .B2(new_n806), .ZN(G1342gat));
  NAND2_X1  g606(.A1(new_n589), .A2(new_n395), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(G134gat), .A3(new_n497), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n797), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n795), .B2(new_n590), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1343gat));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n439), .A3(new_n495), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n466), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n563), .A2(G141gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n693), .A2(new_n793), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n643), .A2(new_n563), .ZN(new_n819));
  INV_X1    g618(.A(new_n788), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n642), .A2(new_n787), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n563), .B2(new_n783), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(new_n590), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n823), .B2(new_n617), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n824), .B2(new_n439), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827), .B2(new_n563), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n817), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n831));
  INV_X1    g630(.A(new_n818), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n791), .B2(new_n441), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n824), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n831), .A2(new_n838), .A3(new_n707), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n839), .A2(G141gat), .B1(new_n815), .B2(new_n816), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n830), .B1(new_n840), .B2(new_n829), .ZN(G1344gat));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n216), .A2(KEYINPUT59), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n831), .A2(new_n838), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n664), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n815), .A2(new_n216), .A3(new_n642), .ZN(new_n846));
  INV_X1    g645(.A(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n834), .A2(new_n835), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n837), .B1(new_n848), .B2(new_n818), .ZN(new_n849));
  AOI211_X1 g648(.A(KEYINPUT118), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n851), .B2(new_n642), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n216), .B1(new_n836), .B2(new_n642), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT119), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n845), .B(new_n846), .C1(new_n852), .C2(new_n855), .ZN(G1345gat));
  AOI21_X1  g655(.A(G155gat), .B1(new_n815), .B2(new_n617), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n617), .A2(G155gat), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT120), .Z(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n851), .B2(new_n859), .ZN(G1346gat));
  OAI21_X1  g659(.A(G162gat), .B1(new_n844), .B2(new_n590), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n808), .A2(G162gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n814), .B2(new_n862), .ZN(G1347gat));
  NOR4_X1   g662(.A1(new_n791), .A2(new_n646), .A3(new_n395), .A4(new_n497), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n328), .A3(new_n707), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n657), .A2(new_n646), .A3(new_n395), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n792), .A2(new_n707), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(KEYINPUT121), .A3(G169gat), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT121), .B1(new_n867), .B2(G169gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1348gat));
  NAND2_X1  g671(.A1(new_n792), .A2(new_n866), .ZN(new_n873));
  OAI21_X1  g672(.A(G176gat), .B1(new_n873), .B2(new_n664), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n329), .A3(new_n642), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1349gat));
  OAI21_X1  g675(.A(G183gat), .B1(new_n873), .B2(new_n663), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n864), .A2(new_n350), .A3(new_n617), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g679(.A(G190gat), .B1(new_n873), .B2(new_n590), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT61), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n334), .A3(new_n589), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1351gat));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n825), .B2(new_n826), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n834), .A2(new_n886), .A3(new_n835), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n646), .A2(new_n395), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n495), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n885), .A2(new_n887), .A3(new_n707), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G197gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n791), .A2(new_n646), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n693), .A2(new_n441), .A3(new_n395), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n310), .A3(new_n707), .A4(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n892), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n893), .A2(new_n894), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(G204gat), .A3(new_n664), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT62), .ZN(new_n904));
  AND4_X1   g703(.A1(new_n642), .A2(new_n885), .A3(new_n887), .A4(new_n890), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n311), .B2(new_n905), .ZN(G1353gat));
  NOR2_X1   g705(.A1(new_n889), .A2(new_n663), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n848), .A2(KEYINPUT126), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(G211gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n848), .A2(new_n907), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AND4_X1   g712(.A1(KEYINPUT63), .A2(new_n912), .A3(G211gat), .A4(new_n908), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n617), .A2(new_n307), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(new_n914), .B1(new_n902), .B2(new_n915), .ZN(G1354gat));
  OAI21_X1  g715(.A(new_n293), .B1(new_n902), .B2(new_n590), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n885), .A2(new_n887), .A3(new_n890), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n589), .A2(G218gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1355gat));
endmodule


