

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n634), .A2(n525), .ZN(n646) );
  AND2_X2 U555 ( .A1(n535), .A2(G2104), .ZN(n885) );
  XNOR2_X1 U556 ( .A(n685), .B(KEYINPUT89), .ZN(n686) );
  INV_X1 U557 ( .A(KEYINPUT91), .ZN(n728) );
  INV_X1 U558 ( .A(KEYINPUT30), .ZN(n685) );
  INV_X1 U559 ( .A(n730), .ZN(n701) );
  XNOR2_X1 U560 ( .A(n687), .B(n686), .ZN(n688) );
  INV_X1 U561 ( .A(KEYINPUT90), .ZN(n726) );
  NOR2_X1 U562 ( .A1(G651), .A2(n634), .ZN(n649) );
  XOR2_X1 U563 ( .A(KEYINPUT68), .B(n577), .Z(n948) );
  NOR2_X1 U564 ( .A1(n543), .A2(n542), .ZN(G160) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U566 ( .A1(n645), .A2(G89), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n521), .B(KEYINPUT4), .ZN(n523) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  INV_X1 U569 ( .A(G651), .ZN(n525) );
  NAND2_X1 U570 ( .A1(G76), .A2(n646), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n524), .B(KEYINPUT5), .ZN(n531) );
  NAND2_X1 U573 ( .A1(G51), .A2(n649), .ZN(n528) );
  NOR2_X1 U574 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X2 U575 ( .A(KEYINPUT1), .B(n526), .Z(n644) );
  NAND2_X1 U576 ( .A1(G63), .A2(n644), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U580 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U581 ( .A(G168), .B(KEYINPUT8), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT71), .ZN(G286) );
  INV_X1 U583 ( .A(G2105), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n885), .A2(G101), .ZN(n534) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n534), .Z(n537) );
  NOR2_X2 U586 ( .A1(G2104), .A2(n535), .ZN(n880) );
  NAND2_X1 U587 ( .A1(n880), .A2(G125), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n538), .B(KEYINPUT64), .ZN(n543) );
  NOR2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT17), .B(n539), .Z(n884) );
  NAND2_X1 U592 ( .A1(G137), .A2(n884), .ZN(n541) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U594 ( .A1(G113), .A2(n881), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G85), .A2(n645), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G72), .A2(n646), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G47), .A2(n649), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G60), .A2(n644), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G290) );
  NAND2_X1 U603 ( .A1(G52), .A2(n649), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G64), .A2(n644), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n646), .A2(G77), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT65), .B(n552), .Z(n554) );
  NAND2_X1 U608 ( .A1(n645), .A2(G90), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U611 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U612 ( .A(G171), .ZN(G301) );
  XOR2_X1 U613 ( .A(G2430), .B(G2443), .Z(n559) );
  XNOR2_X1 U614 ( .A(KEYINPUT95), .B(G2451), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n559), .B(n558), .ZN(n566) );
  XOR2_X1 U616 ( .A(G2435), .B(G2427), .Z(n561) );
  XNOR2_X1 U617 ( .A(G2446), .B(G2454), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U619 ( .A(n562), .B(G2438), .Z(n564) );
  XNOR2_X1 U620 ( .A(G1341), .B(G1348), .ZN(n563) );
  XNOR2_X1 U621 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n566), .B(n565), .ZN(n567) );
  AND2_X1 U623 ( .A1(n567), .A2(G14), .ZN(G401) );
  INV_X1 U624 ( .A(G860), .ZN(n608) );
  NAND2_X1 U625 ( .A1(G68), .A2(n646), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n645), .A2(G81), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n568), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U629 ( .A(n571), .B(KEYINPUT13), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G43), .A2(n649), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n644), .A2(G56), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n574), .Z(n575) );
  NOR2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U635 ( .A1(n608), .A2(n948), .ZN(G153) );
  INV_X1 U636 ( .A(G132), .ZN(G219) );
  INV_X1 U637 ( .A(G82), .ZN(G220) );
  INV_X1 U638 ( .A(G57), .ZN(G237) );
  INV_X1 U639 ( .A(G108), .ZN(G238) );
  INV_X1 U640 ( .A(G120), .ZN(G236) );
  NAND2_X1 U641 ( .A1(n884), .A2(G138), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G126), .A2(n880), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT81), .B(n578), .Z(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G102), .A2(n885), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G114), .A2(n881), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(G164) );
  NAND2_X1 U649 ( .A1(G94), .A2(G452), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT66), .B(n585), .Z(G173) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U653 ( .A(G223), .ZN(n824) );
  NAND2_X1 U654 ( .A1(n824), .A2(G567), .ZN(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G79), .A2(n646), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G54), .A2(n649), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U660 ( .A(KEYINPUT70), .B(n590), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G92), .A2(n645), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G66), .A2(n644), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT69), .B(n593), .Z(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT15), .B(n596), .ZN(n945) );
  INV_X1 U667 ( .A(G868), .ZN(n605) );
  NAND2_X1 U668 ( .A1(n945), .A2(n605), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G53), .A2(n649), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G65), .A2(n644), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G91), .A2(n645), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G78), .A2(n646), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n956) );
  XNOR2_X1 U677 ( .A(n956), .B(KEYINPUT67), .ZN(G299) );
  NAND2_X1 U678 ( .A1(G286), .A2(G868), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G299), .A2(n605), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n608), .A2(G559), .ZN(n609) );
  INV_X1 U682 ( .A(n945), .ZN(n663) );
  NAND2_X1 U683 ( .A1(n609), .A2(n663), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(n948), .A2(G868), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n663), .A2(G868), .ZN(n611) );
  NOR2_X1 U687 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G282) );
  XOR2_X1 U689 ( .A(G2100), .B(KEYINPUT72), .Z(n622) );
  NAND2_X1 U690 ( .A1(n880), .A2(G123), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G111), .A2(n881), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G135), .A2(n884), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G99), .A2(n885), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n988) );
  XNOR2_X1 U698 ( .A(n988), .B(G2096), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U700 ( .A1(G86), .A2(n645), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G48), .A2(n649), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n646), .A2(G73), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n644), .A2(G61), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n649), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U711 ( .A(KEYINPUT76), .B(n632), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n644), .A2(n633), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G88), .A2(n645), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G75), .A2(n646), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G50), .A2(n649), .ZN(n639) );
  XNOR2_X1 U719 ( .A(KEYINPUT77), .B(n639), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(G62), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G67), .A2(n644), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G93), .A2(n645), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G80), .A2(n646), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n649), .A2(G55), .ZN(n650) );
  XOR2_X1 U729 ( .A(KEYINPUT74), .B(n650), .Z(n651) );
  NOR2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n655), .B(KEYINPUT75), .ZN(n837) );
  NOR2_X1 U733 ( .A1(G868), .A2(n837), .ZN(n656) );
  XOR2_X1 U734 ( .A(n656), .B(KEYINPUT78), .Z(n667) );
  XNOR2_X1 U735 ( .A(n837), .B(G288), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(G290), .Z(n657) );
  XNOR2_X1 U737 ( .A(G299), .B(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U739 ( .A(G305), .B(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n948), .B(G166), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n904) );
  NAND2_X1 U742 ( .A1(G559), .A2(n663), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT73), .B(n664), .Z(n834) );
  XNOR2_X1 U744 ( .A(n904), .B(n834), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G236), .A2(G238), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G69), .A2(n672), .ZN(n673) );
  NOR2_X1 U755 ( .A1(n673), .A2(G237), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT79), .ZN(n832) );
  NAND2_X1 U757 ( .A1(n832), .A2(G567), .ZN(n679) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U760 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G96), .A2(n677), .ZN(n831) );
  NAND2_X1 U762 ( .A1(n831), .A2(G2106), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n838), .A2(n680), .ZN(n828) );
  NAND2_X1 U766 ( .A1(n828), .A2(G36), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT80), .B(n681), .ZN(G176) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U769 ( .A(n774), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NAND2_X1 U771 ( .A1(n682), .A2(n775), .ZN(n730) );
  NAND2_X1 U772 ( .A1(G8), .A2(n730), .ZN(n769) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n769), .ZN(n741) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n730), .ZN(n738) );
  INV_X1 U775 ( .A(n738), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G8), .A2(n683), .ZN(n684) );
  OR2_X1 U777 ( .A1(n741), .A2(n684), .ZN(n687) );
  NOR2_X1 U778 ( .A1(G168), .A2(n688), .ZN(n692) );
  XNOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .ZN(n1006) );
  NOR2_X1 U780 ( .A1(n730), .A2(n1006), .ZN(n690) );
  XOR2_X1 U781 ( .A(KEYINPUT86), .B(G1961), .Z(n926) );
  NOR2_X1 U782 ( .A1(n701), .A2(n926), .ZN(n689) );
  NOR2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n721) );
  NOR2_X1 U784 ( .A1(G171), .A2(n721), .ZN(n691) );
  NOR2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n693), .B(KEYINPUT31), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n701), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  INV_X1 U789 ( .A(G1956), .ZN(n957) );
  NOR2_X1 U790 ( .A1(n957), .A2(n701), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n956), .A2(n699), .ZN(n698) );
  XNOR2_X1 U793 ( .A(KEYINPUT28), .B(KEYINPUT87), .ZN(n697) );
  XNOR2_X1 U794 ( .A(n698), .B(n697), .ZN(n719) );
  NAND2_X1 U795 ( .A1(n956), .A2(n699), .ZN(n717) );
  XNOR2_X1 U796 ( .A(KEYINPUT26), .B(KEYINPUT88), .ZN(n707) );
  NOR2_X1 U797 ( .A1(G1996), .A2(n707), .ZN(n700) );
  NOR2_X1 U798 ( .A1(n948), .A2(n700), .ZN(n705) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n730), .ZN(n703) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n701), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n945), .A2(n713), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n712) );
  INV_X1 U804 ( .A(G1341), .ZN(n917) );
  NAND2_X1 U805 ( .A1(n917), .A2(n707), .ZN(n706) );
  NAND2_X1 U806 ( .A1(n706), .A2(n730), .ZN(n710) );
  INV_X1 U807 ( .A(G1996), .ZN(n1007) );
  NOR2_X1 U808 ( .A1(n1007), .A2(n730), .ZN(n708) );
  NAND2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n713), .A2(n945), .ZN(n714) );
  NOR2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U816 ( .A(n720), .B(KEYINPUT29), .ZN(n723) );
  AND2_X1 U817 ( .A1(G171), .A2(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n739) );
  NAND2_X1 U821 ( .A1(n739), .A2(G286), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(n728), .ZN(n735) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n769), .ZN(n732) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U826 ( .A1(G303), .A2(n733), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n736), .A2(G8), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT32), .ZN(n761) );
  NAND2_X1 U830 ( .A1(G8), .A2(n738), .ZN(n743) );
  INV_X1 U831 ( .A(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n762) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n959) );
  AND2_X1 U835 ( .A1(n762), .A2(n959), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n748), .A2(KEYINPUT33), .ZN(n744) );
  OR2_X1 U838 ( .A1(n769), .A2(n744), .ZN(n755) );
  AND2_X1 U839 ( .A1(n745), .A2(n755), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n761), .A2(n746), .ZN(n757) );
  INV_X1 U841 ( .A(n769), .ZN(n752) );
  INV_X1 U842 ( .A(n959), .ZN(n750) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n960) );
  XNOR2_X1 U845 ( .A(KEYINPUT92), .B(n960), .ZN(n749) );
  NOR2_X1 U846 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n753) );
  OR2_X1 U848 ( .A1(KEYINPUT33), .A2(n753), .ZN(n754) );
  NAND2_X1 U849 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U850 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U851 ( .A(G1981), .B(KEYINPUT93), .ZN(n758) );
  XNOR2_X1 U852 ( .A(n758), .B(G305), .ZN(n953) );
  NAND2_X1 U853 ( .A1(n759), .A2(n953), .ZN(n760) );
  XNOR2_X1 U854 ( .A(n760), .B(KEYINPUT94), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n765) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U857 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  AND2_X1 U859 ( .A1(n766), .A2(n769), .ZN(n771) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U861 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  NOR2_X1 U862 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  AND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n807) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n819) );
  NAND2_X1 U866 ( .A1(G140), .A2(n884), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G104), .A2(n885), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(n778), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n880), .A2(G128), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT82), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G116), .A2(n881), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U874 ( .A(n782), .B(KEYINPUT35), .Z(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT36), .B(n785), .Z(n786) );
  XNOR2_X1 U877 ( .A(KEYINPUT83), .B(n786), .ZN(n900) );
  XNOR2_X1 U878 ( .A(KEYINPUT37), .B(G2067), .ZN(n817) );
  NOR2_X1 U879 ( .A1(n900), .A2(n817), .ZN(n996) );
  NAND2_X1 U880 ( .A1(n819), .A2(n996), .ZN(n815) );
  INV_X1 U881 ( .A(n815), .ZN(n804) );
  NAND2_X1 U882 ( .A1(G141), .A2(n884), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G117), .A2(n881), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n885), .A2(G105), .ZN(n789) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n789), .Z(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n880), .A2(G129), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n879) );
  AND2_X1 U890 ( .A1(n879), .A2(G1996), .ZN(n801) );
  NAND2_X1 U891 ( .A1(G131), .A2(n884), .ZN(n795) );
  NAND2_X1 U892 ( .A1(G107), .A2(n881), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U894 ( .A1(G119), .A2(n880), .ZN(n797) );
  NAND2_X1 U895 ( .A1(G95), .A2(n885), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n899) );
  INV_X1 U898 ( .A(G1991), .ZN(n1004) );
  NOR2_X1 U899 ( .A1(n899), .A2(n1004), .ZN(n800) );
  NOR2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n990) );
  INV_X1 U901 ( .A(n819), .ZN(n802) );
  NOR2_X1 U902 ( .A1(n990), .A2(n802), .ZN(n812) );
  XNOR2_X1 U903 ( .A(KEYINPUT84), .B(n812), .ZN(n803) );
  NOR2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U905 ( .A(n805), .B(KEYINPUT85), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n947) );
  NAND2_X1 U908 ( .A1(n947), .A2(n819), .ZN(n808) );
  NAND2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n822) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n879), .ZN(n982) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n810) );
  AND2_X1 U912 ( .A1(n1004), .A2(n899), .ZN(n992) );
  NOR2_X1 U913 ( .A1(n810), .A2(n992), .ZN(n811) );
  NOR2_X1 U914 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U915 ( .A1(n982), .A2(n813), .ZN(n814) );
  XNOR2_X1 U916 ( .A(n814), .B(KEYINPUT39), .ZN(n816) );
  NAND2_X1 U917 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U918 ( .A1(n900), .A2(n817), .ZN(n997) );
  NAND2_X1 U919 ( .A1(n818), .A2(n997), .ZN(n820) );
  NAND2_X1 U920 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U921 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n823), .ZN(G329) );
  NAND2_X1 U923 ( .A1(n824), .A2(G2106), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n825), .B(KEYINPUT96), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n826) );
  XNOR2_X1 U926 ( .A(KEYINPUT97), .B(n826), .ZN(n827) );
  NAND2_X1 U927 ( .A1(n827), .A2(G661), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U929 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n830), .B(KEYINPUT98), .ZN(G188) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n833), .B(KEYINPUT99), .ZN(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U936 ( .A(n948), .B(n834), .ZN(n835) );
  NOR2_X1 U937 ( .A1(G860), .A2(n835), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(G145) );
  INV_X1 U939 ( .A(n838), .ZN(G319) );
  XOR2_X1 U940 ( .A(KEYINPUT103), .B(G1976), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1956), .B(G1981), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G1971), .B(G1961), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1966), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT102), .B(G2474), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U953 ( .A(KEYINPUT100), .B(G2678), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U958 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2100), .B(G2096), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n880), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n860), .B(KEYINPUT44), .ZN(n861) );
  XNOR2_X1 U965 ( .A(KEYINPUT104), .B(n861), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G100), .A2(n885), .ZN(n862) );
  XOR2_X1 U967 ( .A(KEYINPUT105), .B(n862), .Z(n863) );
  NAND2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G136), .A2(n884), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G112), .A2(n881), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U972 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  NAND2_X1 U974 ( .A1(G139), .A2(n884), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G103), .A2(n885), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G127), .A2(n880), .ZN(n872) );
  NAND2_X1 U978 ( .A1(G115), .A2(n881), .ZN(n871) );
  NAND2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U980 ( .A(KEYINPUT47), .B(n873), .ZN(n874) );
  XNOR2_X1 U981 ( .A(KEYINPUT107), .B(n874), .ZN(n875) );
  NOR2_X1 U982 ( .A1(n876), .A2(n875), .ZN(n975) );
  XNOR2_X1 U983 ( .A(n975), .B(KEYINPUT108), .ZN(n877) );
  XNOR2_X1 U984 ( .A(n878), .B(n877), .ZN(n898) );
  XOR2_X1 U985 ( .A(n879), .B(G162), .Z(n893) );
  NAND2_X1 U986 ( .A1(G130), .A2(n880), .ZN(n883) );
  NAND2_X1 U987 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U988 ( .A1(n883), .A2(n882), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G142), .A2(n884), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G106), .A2(n885), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(KEYINPUT106), .B(n888), .Z(n889) );
  XNOR2_X1 U993 ( .A(KEYINPUT45), .B(n889), .ZN(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n988), .B(n894), .Z(n896) );
  XNOR2_X1 U997 ( .A(G164), .B(G160), .ZN(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT109), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n945), .B(G286), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(G301), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT110), .B(n909), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(KEYINPUT111), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n911), .B(n910), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n912), .B(KEYINPUT112), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n915), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n916), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1019 ( .A(G19), .B(n917), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G1956), .B(G20), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1025 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT60), .B(n925), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n926), .B(G5), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G21), .B(G1966), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(KEYINPUT122), .B(n931), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n938) );
  XNOR2_X1 U1034 ( .A(G1986), .B(G24), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G1971), .B(KEYINPUT123), .ZN(n934) );
  XNOR2_X1 U1038 ( .A(n934), .B(G22), .ZN(n935) );
  NAND2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1040 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n941), .B(KEYINPUT61), .ZN(n942) );
  XOR2_X1 U1043 ( .A(KEYINPUT125), .B(n942), .Z(n943) );
  NOR2_X1 U1044 ( .A1(G16), .A2(n943), .ZN(n973) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT119), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(n944), .B(KEYINPUT56), .ZN(n971) );
  XNOR2_X1 U1047 ( .A(G1348), .B(n945), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G301), .B(G1961), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G1341), .B(n948), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n969) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(n955), .B(KEYINPUT57), .ZN(n967) );
  NAND2_X1 U1056 ( .A1(G303), .A2(G1971), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n956), .B(KEYINPUT120), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(n958), .B(n957), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(KEYINPUT121), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT126), .ZN(n1003) );
  XNOR2_X1 U1068 ( .A(G164), .B(G2078), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G2072), .B(n975), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT114), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT50), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT115), .B(n980), .Z(n985) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(KEYINPUT51), .B(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(G160), .B(G2084), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT113), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n999), .ZN(n1000) );
  OR2_X1 U1087 ( .A1(KEYINPUT55), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1029) );
  XOR2_X1 U1090 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n1024) );
  XNOR2_X1 U1091 ( .A(G2090), .B(G35), .ZN(n1019) );
  XNOR2_X1 U1092 ( .A(G25), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(G28), .ZN(n1016) );
  XOR2_X1 U1094 ( .A(n1006), .B(G27), .Z(n1009) );
  XOR2_X1 U1095 ( .A(n1007), .B(G32), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT116), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G2067), .B(G26), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G33), .B(G2072), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1105 ( .A(G2084), .B(G34), .Z(n1020) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1024), .B(n1023), .ZN(n1025) );
  OR2_X1 U1109 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(G11), .A2(n1026), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT118), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(n1030), .B(KEYINPUT62), .Z(n1031) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1031), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

