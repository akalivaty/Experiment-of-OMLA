//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT77), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  AOI21_X1  g0051(.A(G1), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G274), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n252), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT65), .B(G226), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n261), .B1(new_n224), .B2(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AOI211_X1 g0064(.A(new_n254), .B(new_n258), .C1(new_n264), .C2(new_n255), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n205), .A2(KEYINPUT66), .A3(G20), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT66), .B1(new_n205), .B2(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n214), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(G50), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n206), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G58), .A2(G68), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n206), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n277), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n275), .A2(new_n287), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n279), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT9), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n265), .A2(G190), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n267), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n267), .A2(new_n292), .A3(new_n296), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n265), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n291), .B1(new_n265), .B2(G169), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n278), .A2(G68), .A3(new_n271), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n275), .A2(new_n218), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT12), .ZN(new_n306));
  INV_X1    g0106(.A(new_n277), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n206), .A2(G33), .A3(G77), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT11), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n259), .A2(G226), .A3(new_n260), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G97), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(new_n248), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n255), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n254), .B1(G238), .B2(new_n256), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(new_n321), .A3(new_n320), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G190), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n322), .A2(new_n323), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT14), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n326), .A2(G179), .A3(new_n327), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n314), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G107), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n341), .B1(new_n345), .B2(new_n259), .C1(new_n262), .C2(new_n219), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n255), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n254), .B1(G244), .B2(new_n256), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(KEYINPUT68), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n271), .A2(G77), .A3(new_n278), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G77), .B2(new_n274), .ZN(new_n356));
  INV_X1    g0156(.A(new_n280), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n281), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n307), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n354), .B(new_n363), .C1(new_n266), .C2(new_n353), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n353), .B2(new_n299), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n351), .A2(new_n332), .A3(new_n352), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n302), .A2(new_n340), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n270), .A2(new_n280), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n278), .B1(new_n275), .B2(new_n280), .ZN(new_n372));
  NAND3_X1  g0172(.A1(KEYINPUT71), .A2(G58), .A3(G68), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT71), .B1(G58), .B2(G68), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n374), .A2(new_n375), .A3(new_n286), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n376), .A2(new_n206), .B1(new_n377), .B2(new_n284), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G33), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g0184(.A(G20), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n218), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n384), .ZN(new_n388));
  AND2_X1   g0188(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(G33), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(G20), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n378), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n307), .B1(new_n394), .B2(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n248), .B1(new_n389), .B2(new_n390), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n380), .A2(G33), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n384), .A2(new_n398), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n400), .B2(new_n206), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n375), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n373), .C1(G58), .C2(G68), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT73), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n410), .B(new_n407), .C1(new_n402), .C2(new_n405), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n395), .B(KEYINPUT74), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n386), .B1(new_n259), .B2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(new_n398), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n248), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n417), .B2(new_n396), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n378), .B1(new_n418), .B2(G68), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n410), .B1(new_n419), .B2(new_n407), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n406), .A2(KEYINPUT73), .A3(new_n408), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT74), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n372), .B1(new_n413), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n256), .A2(G232), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n253), .ZN(new_n426));
  MUX2_X1   g0226(.A(G223), .B(G226), .S(G1698), .Z(new_n427));
  NAND2_X1  g0227(.A1(new_n392), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n430), .B2(new_n255), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G179), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n250), .B1(new_n428), .B2(new_n429), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT75), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n432), .B2(new_n434), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n424), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT18), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n431), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(new_n446), .C1(G200), .C2(new_n431), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n372), .B(new_n447), .C1(new_n413), .C2(new_n423), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n372), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n395), .B1(new_n409), .B2(new_n411), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n454), .B2(new_n412), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n447), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n424), .A2(new_n457), .A3(new_n439), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n441), .A2(new_n450), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n247), .B1(new_n370), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n459), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(KEYINPUT77), .A3(new_n369), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G33), .B1(new_n381), .B2(new_n382), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT7), .B(new_n206), .C1(new_n465), .C2(new_n415), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n345), .B1(new_n466), .B2(new_n414), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n468), .A2(new_n317), .A3(G107), .ZN(new_n469));
  XNOR2_X1  g0269(.A(G97), .B(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n471), .A2(new_n206), .B1(new_n224), .B2(new_n284), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n277), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n275), .A2(new_n317), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n205), .A2(G33), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n307), .A2(new_n274), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n476), .B2(new_n317), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT78), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G33), .A3(G283), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n383), .A2(new_n384), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n225), .A2(G1698), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n250), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G274), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n255), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT80), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n249), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(G41), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT79), .A3(new_n205), .A4(G45), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n205), .B(G45), .C1(new_n249), .C2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n495), .A2(new_n501), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(G41), .B1(new_n497), .B2(new_n499), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(new_n250), .C1(new_n508), .C2(new_n504), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n332), .B1(new_n493), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT4), .B1(new_n392), .B2(new_n490), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n255), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(KEYINPUT81), .A3(new_n509), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n516), .A3(new_n299), .A4(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n479), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT82), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n513), .A2(new_n516), .A3(new_n522), .A4(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(G200), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n507), .A3(new_n509), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n473), .B(new_n478), .C1(new_n525), .C2(new_n442), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT83), .B(G116), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n476), .A2(new_n529), .B1(new_n531), .B2(new_n274), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n206), .B1(new_n317), .B2(G33), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n483), .B2(new_n485), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n530), .A2(G20), .B1(new_n214), .B2(new_n276), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT20), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G270), .B(new_n250), .C1(new_n508), .C2(new_n504), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G257), .A2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n227), .B2(G1698), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n392), .A2(new_n543), .B1(G303), .B2(new_n400), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n507), .B(new_n541), .C1(new_n544), .C2(new_n250), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n540), .A2(G169), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n539), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n537), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n532), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n392), .A2(new_n543), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n400), .A2(G303), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n250), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n507), .A2(new_n541), .ZN(new_n555));
  OAI21_X1  g0355(.A(G200), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n556), .C1(new_n442), .C2(new_n545), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n545), .A2(new_n299), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n540), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT21), .A4(G169), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n548), .A2(new_n557), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n221), .B1(new_n251), .B2(G1), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n205), .A2(new_n494), .A3(G45), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n250), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n225), .B2(G1698), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n383), .A3(new_n384), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n531), .A2(G33), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n565), .B1(new_n570), .B2(new_n250), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n332), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G87), .A2(G97), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n342), .A2(new_n344), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n206), .B1(new_n248), .B2(new_n317), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n281), .A2(KEYINPUT19), .A3(new_n317), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n206), .A2(G68), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n577), .A2(new_n578), .B1(new_n489), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n277), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n275), .A2(new_n359), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n476), .A2(new_n359), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n250), .B1(new_n568), .B2(new_n569), .ZN(new_n585));
  INV_X1    g0385(.A(new_n565), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n299), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n572), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G190), .B(new_n565), .C1(new_n570), .C2(new_n250), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n580), .A2(new_n277), .B1(new_n275), .B2(new_n359), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n278), .A2(G87), .A3(new_n475), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n528), .A2(new_n562), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n206), .A2(G87), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n400), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n342), .A2(new_n344), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT23), .B1(new_n601), .B2(new_n206), .ZN(new_n602));
  OR3_X1    g0402(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n383), .A2(KEYINPUT22), .A3(G87), .A4(new_n384), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(new_n569), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n604), .B(new_n605), .C1(new_n607), .C2(G20), .ZN(new_n608));
  AOI21_X1  g0408(.A(G20), .B1(new_n606), .B2(new_n569), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT24), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n277), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT25), .B1(new_n275), .B2(new_n226), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n226), .B2(new_n476), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(G264), .B(new_n250), .C1(new_n508), .C2(new_n504), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n221), .A2(new_n260), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n260), .A2(G257), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n383), .A2(new_n384), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(G33), .A2(G294), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n250), .B1(new_n626), .B2(KEYINPUT84), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n507), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n332), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n299), .A3(new_n507), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n619), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n617), .B1(new_n612), .B2(new_n277), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n630), .A2(new_n442), .A3(new_n507), .ZN(new_n636));
  AOI21_X1  g0436(.A(G200), .B1(new_n630), .B2(new_n507), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n634), .A2(KEYINPUT85), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT85), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n597), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n464), .A2(new_n641), .ZN(G372));
  NOR2_X1   g0442(.A1(new_n300), .A2(new_n301), .ZN(new_n643));
  INV_X1    g0443(.A(new_n435), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT18), .B1(new_n455), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n424), .A2(new_n457), .A3(new_n435), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n367), .A2(new_n330), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n338), .B2(new_n337), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n450), .A2(new_n456), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n645), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n650), .A2(new_n651), .B1(new_n295), .B2(new_n297), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n643), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n565), .A2(KEYINPUT86), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT86), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n250), .A2(new_n563), .A3(new_n564), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(G200), .B1(new_n585), .B2(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n591), .A2(new_n590), .A3(new_n593), .A4(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n332), .B1(new_n585), .B2(new_n658), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT87), .B(new_n332), .C1(new_n585), .C2(new_n658), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n584), .A3(new_n588), .A4(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n519), .A2(new_n661), .A3(new_n662), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n479), .A2(new_n511), .A3(new_n518), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT26), .B1(new_n595), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n672), .A2(new_n671), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT90), .A3(new_n668), .A4(new_n670), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n527), .A2(new_n524), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n665), .A2(new_n666), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n584), .A2(new_n588), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n660), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n679), .A2(new_n638), .A3(new_n682), .A4(new_n669), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n528), .A2(KEYINPUT88), .A3(new_n638), .A4(new_n682), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n548), .A2(new_n560), .A3(new_n559), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n634), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n654), .B1(new_n464), .B2(new_n691), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n273), .A2(new_n206), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(G213), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n639), .A2(new_n640), .B1(new_n635), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n702), .B(new_n703), .C1(new_n634), .C2(new_n699), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n687), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n551), .A2(new_n699), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n561), .B2(new_n707), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n702), .A2(new_n703), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n687), .A2(new_n698), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n634), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n699), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n209), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n575), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n212), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n597), .B(new_n699), .C1(new_n640), .C2(new_n639), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n493), .A2(new_n510), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n558), .A2(new_n731), .A3(new_n587), .ZN(new_n732));
  INV_X1    g0532(.A(new_n630), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n525), .A2(new_n571), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n630), .A4(new_n558), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n585), .A2(new_n658), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(new_n545), .A3(new_n299), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n631), .A3(new_n520), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n740), .B2(new_n698), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n711), .B1(new_n729), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n682), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT26), .B1(new_n745), .B2(new_n669), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n596), .A2(new_n662), .A3(new_n519), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n676), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n687), .A2(new_n634), .ZN(new_n749));
  OR3_X1    g0549(.A1(new_n749), .A2(new_n683), .A3(KEYINPUT93), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT93), .B1(new_n749), .B2(new_n683), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n698), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n690), .A2(new_n699), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n744), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n728), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n272), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n205), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n723), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n712), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n710), .A2(new_n711), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n710), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n214), .B1(G20), .B2(new_n332), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n206), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n220), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n442), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n400), .B(new_n774), .C1(G107), .C2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT95), .Z(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G159), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(new_n299), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n442), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n779), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G68), .B1(new_n788), .B2(G77), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n299), .A2(new_n266), .A3(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n317), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n266), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G58), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n287), .A2(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n793), .B(new_n800), .C1(KEYINPUT32), .C2(new_n782), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n778), .A2(new_n783), .A3(new_n789), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n798), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G294), .B2(new_n791), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n400), .B1(new_n773), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT96), .Z(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n785), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n812), .A2(new_n775), .B1(new_n787), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n814), .C1(G329), .C2(new_n781), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n806), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n771), .B1(new_n802), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n763), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n768), .A2(new_n770), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n722), .A2(new_n392), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n251), .B2(new_n213), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n242), .A2(new_n251), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n209), .A2(new_n259), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n825), .A2(new_n203), .B1(G116), .B2(new_n209), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n823), .A2(new_n824), .B1(KEYINPUT94), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(KEYINPUT94), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n820), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n817), .A2(new_n818), .A3(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n764), .A2(new_n765), .B1(new_n769), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n368), .A2(new_n698), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n690), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n755), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n367), .A2(new_n698), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n364), .B1(new_n363), .B2(new_n699), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n367), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n744), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n763), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n770), .A2(new_n766), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n763), .B1(G77), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT97), .Z(new_n847));
  NOR2_X1   g0647(.A1(new_n775), .A2(new_n218), .ZN(new_n848));
  INV_X1    g0648(.A(new_n773), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G50), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n780), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n489), .B(new_n852), .C1(G58), .C2(new_n791), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n786), .A2(G150), .B1(new_n788), .B2(G159), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(new_n798), .B2(new_n855), .C1(new_n856), .C2(new_n796), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT34), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n853), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n793), .B1(G294), .B2(new_n797), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT99), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n400), .B1(new_n775), .B2(new_n220), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n773), .A2(new_n226), .B1(new_n780), .B2(new_n813), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(G303), .C2(new_n795), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n785), .A2(new_n812), .B1(new_n787), .B2(new_n530), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT98), .Z(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n847), .B1(new_n771), .B2(new_n870), .C1(new_n838), .C2(new_n767), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT100), .Z(new_n872));
  NOR2_X1   g0672(.A1(new_n843), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(G384));
  OAI21_X1  g0674(.A(new_n395), .B1(new_n394), .B2(new_n407), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n696), .B1(new_n875), .B2(new_n372), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n459), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n696), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n424), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n440), .A2(new_n879), .A3(new_n880), .A4(new_n448), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n644), .A2(new_n696), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n875), .A2(new_n372), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n448), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n882), .B1(new_n881), .B2(new_n887), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n877), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n448), .B1(new_n455), .B2(new_n696), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n455), .A2(new_n644), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n881), .ZN(new_n894));
  INV_X1    g0694(.A(new_n879), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n645), .A2(new_n646), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n649), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n890), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n877), .B1(new_n888), .B2(new_n889), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n899), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n337), .A2(new_n338), .A3(new_n699), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n314), .A2(new_n699), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n337), .B2(new_n330), .ZN(new_n911));
  INV_X1    g0711(.A(new_n910), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT103), .B1(new_n339), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n336), .A2(new_n334), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n326), .A2(new_n327), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n335), .B1(new_n915), .B2(G169), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n338), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND4_X1   g0717(.A1(KEYINPUT103), .A2(new_n917), .A3(new_n329), .A4(new_n912), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n911), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n365), .A2(new_n366), .A3(new_n699), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT101), .Z(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT102), .B1(new_n834), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n924), .B(new_n921), .C1(new_n690), .C2(new_n833), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n905), .A2(new_n890), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(new_n896), .B2(new_n696), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n909), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n463), .A2(new_n754), .A3(new_n757), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n654), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT105), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n930), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n436), .A2(new_n438), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n880), .B1(new_n455), .B2(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n455), .A2(new_n447), .B1(new_n884), .B2(new_n883), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n891), .A2(new_n938), .B1(new_n939), .B2(new_n880), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT104), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n941), .A2(new_n942), .B1(new_n459), .B2(new_n876), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n936), .B1(new_n943), .B2(KEYINPUT38), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n729), .A2(new_n743), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n945), .A2(new_n919), .A3(KEYINPUT40), .A4(new_n838), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n935), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n901), .A2(KEYINPUT106), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n919), .A3(new_n838), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n905), .B2(new_n890), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n950), .B1(KEYINPUT40), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n463), .A2(new_n945), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n934), .A2(new_n956), .B1(new_n205), .B2(new_n760), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n934), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n471), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(G116), .A3(new_n215), .A4(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT36), .Z(new_n963));
  NAND4_X1  g0763(.A1(new_n403), .A2(new_n213), .A3(G77), .A4(new_n373), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n287), .A2(G68), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n205), .B(G13), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n958), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT107), .Z(G367));
  NAND2_X1  g0768(.A1(new_n479), .A2(new_n698), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n528), .A2(new_n969), .B1(new_n519), .B2(new_n698), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n715), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n970), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n718), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT108), .Z(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT109), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n719), .A2(new_n679), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n698), .B1(new_n978), .B2(new_n669), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n975), .B2(KEYINPUT42), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n591), .A2(new_n593), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n676), .A2(new_n983), .A3(new_n699), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n682), .B1(new_n983), .B2(new_n699), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n977), .A2(new_n981), .ZN(new_n989));
  INV_X1    g0789(.A(new_n987), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n989), .A2(new_n971), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n988), .A2(new_n991), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n982), .A2(new_n972), .A3(new_n987), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n971), .B1(new_n989), .B2(new_n990), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n723), .B(KEYINPUT41), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n720), .A2(new_n973), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n720), .A2(new_n973), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n715), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n718), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n704), .B2(new_n717), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n712), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n758), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n997), .B1(new_n1009), .B2(new_n758), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n992), .B(new_n996), .C1(new_n762), .C2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n819), .B1(new_n209), .B2(new_n359), .C1(new_n822), .C2(new_n238), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n763), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT110), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n855), .A2(new_n796), .B1(new_n798), .B2(new_n282), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n792), .A2(new_n218), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n785), .A2(new_n377), .B1(new_n787), .B2(new_n287), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n775), .A2(new_n224), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n259), .B1(new_n773), .B2(new_n799), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G137), .C2(new_n781), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n788), .A2(G283), .B1(new_n601), .B2(new_n791), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT111), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n780), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n775), .A2(new_n317), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G294), .C2(new_n786), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n797), .A2(G303), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n392), .B1(G311), .B2(new_n795), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT46), .B1(new_n773), .B2(new_n529), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n530), .A2(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n773), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1024), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT47), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n770), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n768), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1014), .B1(new_n1039), .B2(new_n1041), .C1(new_n986), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1011), .A2(new_n1043), .ZN(G387));
  OAI22_X1  g0844(.A1(new_n775), .A2(new_n530), .B1(new_n780), .B2(new_n804), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n786), .A2(G311), .B1(new_n788), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n798), .B2(new_n1027), .C1(new_n803), .C2(new_n796), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(G294), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(new_n812), .B2(new_n792), .C1(new_n1050), .C2(new_n773), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n392), .B(new_n1045), .C1(new_n1053), .C2(KEYINPUT49), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(KEYINPUT49), .B2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n792), .A2(new_n359), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n798), .A2(new_n287), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G159), .C2(new_n795), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n788), .A2(G68), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n786), .A2(new_n357), .B1(new_n781), .B2(G150), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n489), .B(new_n1029), .C1(G77), .C2(new_n849), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n771), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n821), .B1(new_n235), .B2(new_n251), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n725), .B2(new_n825), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n280), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT113), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n725), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1065), .A2(new_n1071), .B1(new_n226), .B2(new_n722), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n763), .B1(new_n1072), .B2(new_n820), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1063), .B(new_n1073), .C1(new_n705), .C2(new_n768), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1006), .B2(new_n762), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1007), .A2(new_n723), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1006), .A2(new_n758), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  AOI21_X1  g0878(.A(new_n715), .B1(new_n999), .B2(new_n1001), .ZN(new_n1079));
  MUX2_X1   g0879(.A(new_n1003), .B(new_n1079), .S(KEYINPUT114), .Z(new_n1080));
  OAI211_X1 g0880(.A(new_n723), .B(new_n1009), .C1(new_n1080), .C2(new_n1008), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G150), .A2(new_n795), .B1(new_n797), .B2(G159), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n785), .A2(new_n287), .B1(new_n780), .B2(new_n855), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n357), .B2(new_n788), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n775), .A2(new_n220), .B1(new_n773), .B2(new_n218), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n792), .A2(new_n224), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n489), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(KEYINPUT51), .B2(new_n1083), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G311), .A2(new_n797), .B1(new_n795), .B2(G317), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT116), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G294), .A2(new_n788), .B1(new_n781), .B2(G322), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n812), .B2(new_n773), .C1(new_n807), .C2(new_n785), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n400), .B1(new_n775), .B2(new_n226), .C1(new_n792), .C2(new_n530), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n770), .B1(new_n1091), .B2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n821), .A2(new_n245), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n819), .B1(new_n317), .B2(new_n209), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1100), .B(new_n763), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n970), .B2(new_n768), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1080), .B2(new_n762), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1081), .A2(new_n1105), .ZN(G390));
  OAI22_X1  g0906(.A1(new_n787), .A2(new_n317), .B1(new_n780), .B2(new_n1050), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n848), .B(new_n1107), .C1(new_n601), .C2(new_n786), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n529), .A2(new_n798), .B1(new_n796), .B2(new_n812), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1109), .A2(new_n1088), .A3(new_n259), .A4(new_n774), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n259), .B1(new_n856), .B2(new_n785), .C1(new_n798), .C2(new_n851), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n787), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n775), .A2(new_n287), .B1(new_n780), .B2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n773), .A2(new_n282), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n796), .A2(new_n1120), .B1(new_n377), .B2(new_n792), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1108), .A2(new_n1110), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n763), .B1(new_n357), .B2(new_n845), .C1(new_n1123), .C2(new_n771), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n907), .B2(new_n766), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n744), .A2(new_n838), .A3(new_n919), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(KEYINPUT117), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n903), .A2(new_n906), .B1(new_n926), .B2(new_n908), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n921), .B1(new_n753), .B2(new_n838), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n919), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n908), .B(new_n901), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1129), .B(new_n1130), .C1(new_n1131), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n926), .A2(new_n908), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n907), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1138), .A2(new_n1128), .A3(new_n1127), .A4(new_n1134), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1125), .B1(new_n1140), .B2(new_n762), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n463), .A2(new_n744), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n931), .A2(new_n654), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT118), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n931), .A2(KEYINPUT118), .A3(new_n1142), .A4(new_n654), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n838), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1133), .B1(new_n840), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1126), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n923), .B2(new_n925), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1132), .A2(new_n1126), .A3(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n724), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1136), .A2(new_n1153), .A3(new_n1139), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1136), .A2(new_n1153), .A3(new_n1139), .A4(KEYINPUT119), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1141), .B1(new_n1162), .B2(new_n1163), .ZN(G378));
  NAND2_X1  g0964(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT106), .B1(new_n901), .B2(new_n948), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n935), .B(new_n946), .C1(new_n890), .C2(new_n900), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(G330), .B1(new_n952), .B2(KEYINPUT40), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT122), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n951), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n890), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n941), .A2(new_n942), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT38), .B1(new_n1176), .B2(new_n877), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT40), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n711), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT122), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n950), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n291), .A2(new_n878), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n302), .B(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1173), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT123), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n1186), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1173), .A2(new_n1182), .A3(new_n1189), .A4(new_n1187), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1192), .A2(new_n930), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n930), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1168), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n930), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1180), .A2(new_n950), .A3(new_n1186), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT123), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1180), .A2(new_n950), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1186), .B1(new_n1200), .B2(KEYINPUT122), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1199), .B1(new_n1201), .B2(new_n1182), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1193), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1192), .A2(new_n930), .A3(new_n1193), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1166), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1196), .B(new_n723), .C1(new_n1206), .C2(KEYINPUT57), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1187), .A2(new_n766), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n763), .B1(G50), .B2(new_n845), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n392), .A2(G41), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1211), .C1(new_n248), .C2(new_n249), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G97), .A2(new_n786), .B1(new_n776), .B2(G58), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n1211), .C1(new_n359), .C2(new_n787), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n226), .A2(new_n798), .B1(new_n796), .B2(new_n529), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n773), .A2(new_n224), .B1(new_n780), .B2(new_n812), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1016), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1212), .B1(new_n1217), .B2(KEYINPUT58), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n796), .A2(new_n1114), .B1(new_n282), .B2(new_n792), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n788), .A2(G137), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n851), .B2(new_n785), .C1(new_n773), .C2(new_n1112), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G128), .C2(new_n797), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n248), .B(new_n249), .C1(new_n775), .C2(new_n377), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G124), .B2(new_n781), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT59), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1218), .B1(KEYINPUT58), .B2(new_n1217), .C1(new_n1224), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1210), .B1(new_n1229), .B2(new_n770), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1208), .A2(new_n762), .B1(new_n1209), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1207), .A2(new_n1231), .ZN(G375));
  NAND3_X1  g1032(.A1(new_n1165), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n997), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1153), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n812), .A2(new_n798), .B1(new_n796), .B2(new_n1050), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1236), .A2(new_n1056), .A3(new_n259), .A4(new_n1021), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n785), .A2(new_n530), .B1(new_n773), .B2(new_n317), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n345), .A2(new_n787), .B1(new_n780), .B2(new_n807), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n851), .A2(new_n796), .B1(new_n798), .B2(new_n856), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G50), .B2(new_n791), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n781), .A2(G128), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n282), .B2(new_n787), .C1(new_n785), .C2(new_n1112), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n775), .A2(new_n799), .B1(new_n773), .B2(new_n377), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n489), .A3(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1237), .A2(new_n1240), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n763), .B1(G68), .B2(new_n845), .C1(new_n1247), .C2(new_n771), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1133), .B2(new_n766), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1152), .B2(new_n762), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1235), .A2(new_n1250), .ZN(G381));
  OR4_X1    g1051(.A1(G396), .A2(G393), .A3(G381), .A4(G384), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(G387), .A2(G390), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G375), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1160), .A2(new_n1141), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(G407));
  NAND2_X1  g1057(.A1(new_n697), .A2(G213), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G375), .C2(new_n1260), .ZN(G409));
  XNOR2_X1  g1061(.A(G393), .B(G396), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1081), .A2(new_n1105), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1081), .B2(new_n1105), .ZN(new_n1264));
  OAI21_X1  g1064(.A(G387), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1262), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G390), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1081), .A2(new_n1105), .A3(new_n1262), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1011), .A3(new_n1043), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n723), .B1(new_n1272), .B2(new_n1233), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1233), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1250), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(new_n873), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n873), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1259), .A2(G2897), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1206), .A2(new_n1234), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1255), .B1(new_n1231), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1207), .A2(G378), .A3(new_n1231), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1207), .A2(G378), .A3(KEYINPUT125), .A4(new_n1231), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1287), .B2(new_n1259), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1287), .A2(new_n1259), .A3(new_n1278), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1271), .B(new_n1288), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1282), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1259), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1278), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1270), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(G387), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1267), .A2(new_n1268), .B1(new_n1011), .B2(new_n1043), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1288), .A2(new_n1271), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1289), .A2(KEYINPUT63), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1302), .A2(new_n1303), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n1307), .ZN(G405));
  OAI21_X1  g1108(.A(new_n1292), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1309), .B1(new_n1312), .B2(new_n1310), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1265), .A2(new_n1269), .A3(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1302), .A2(KEYINPUT127), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


