//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n439, new_n450, new_n451, new_n453,
    new_n455, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n466, new_n467, new_n468, new_n469, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  OR2_X1    g012(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(new_n439), .ZN(G220));
  INV_X1    g015(.A(G96), .ZN(G221));
  INV_X1    g016(.A(G69), .ZN(G235));
  INV_X1    g017(.A(G120), .ZN(G236));
  INV_X1    g018(.A(G57), .ZN(G237));
  INV_X1    g019(.A(G108), .ZN(G238));
  NAND4_X1  g020(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  INV_X1    g027(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n453), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n453), .A2(G2106), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G217));
  NOR3_X1   g031(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n438), .A2(new_n439), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR4_X1   g036(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g039(.A(G261), .ZN(G325));
  NAND2_X1  g040(.A1(new_n460), .A2(G2106), .ZN(new_n466));
  INV_X1    g041(.A(G567), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G319));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n479), .A2(G137), .B1(G101), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n478), .A2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n479), .A2(G136), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n480), .B1(new_n475), .B2(new_n476), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n491), .B(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n494), .B2(new_n495), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n503), .B(new_n506), .C1(new_n495), .C2(new_n494), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(G50), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n515), .A2(KEYINPUT73), .A3(G50), .A4(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(G75), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(G651), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n511), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n520), .A2(new_n521), .B1(new_n525), .B2(new_n509), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n524), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND2_X1  g104(.A1(new_n515), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT75), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n525), .B2(new_n509), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n526), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n520), .A2(new_n521), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n541), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n537), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n541), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n536), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n526), .A2(G90), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(new_n521), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n519), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n546), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n536), .A2(G43), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT77), .B(G81), .Z(new_n560));
  NAND2_X1  g135(.A1(new_n526), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n520), .B2(new_n521), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT79), .B(new_n573), .C1(new_n553), .C2(new_n571), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(G651), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n533), .A2(new_n580), .A3(G53), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n579), .A2(new_n581), .B1(G91), .B2(new_n526), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  NAND3_X1  g158(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n526), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n541), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n533), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n526), .A2(G86), .B1(new_n533), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n541), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT80), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n546), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI211_X1 g171(.A(KEYINPUT81), .B(new_n546), .C1(new_n591), .C2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n546), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n536), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(new_n526), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n526), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n541), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n546), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n536), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G860), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n611), .B1(G559), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT83), .Z(G148));
  NOR2_X1   g197(.A1(new_n611), .A2(G559), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g202(.A(KEYINPUT3), .B(G2104), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n481), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n479), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n489), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n480), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT86), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT87), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT88), .Z(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n677), .A2(new_n682), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n693), .B1(new_n691), .B2(new_n694), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n674), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n673), .A3(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  NOR2_X1   g277(.A1(G29), .A2(G35), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G162), .B2(G29), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT29), .Z(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT103), .ZN(new_n708));
  NOR2_X1   g283(.A1(G4), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n612), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT95), .B(G1348), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  INV_X1    g287(.A(G1341), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n562), .A2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G19), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n712), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G26), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n489), .A2(G128), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G140), .ZN(new_n723));
  OR2_X1    g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n719), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2067), .ZN(new_n729));
  INV_X1    g304(.A(new_n717), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G1341), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n718), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n718), .A2(KEYINPUT96), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n708), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n719), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n489), .A2(G129), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT99), .Z(new_n739));
  AND2_X1   g314(.A1(new_n481), .A2(G105), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n740), .B(new_n742), .C1(G141), .C2(new_n479), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT100), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g324(.A1(G301), .A2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n715), .A2(G5), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  NAND2_X1  g329(.A1(G160), .A2(G29), .ZN(new_n755));
  AND2_X1   g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NOR2_X1   g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n719), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT98), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n746), .B2(new_n747), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT102), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n749), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n766));
  NAND2_X1  g341(.A1(G103), .A2(G2104), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G2105), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n480), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n479), .A2(G139), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n480), .B2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G33), .B(new_n772), .S(G29), .Z(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2072), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(KEYINPUT97), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(KEYINPUT97), .ZN(new_n777));
  INV_X1    g352(.A(G1966), .ZN(new_n778));
  NOR2_X1   g353(.A1(G168), .A2(new_n715), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n715), .B2(G21), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n773), .A2(G2072), .ZN(new_n783));
  NOR2_X1   g358(.A1(G27), .A2(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G164), .B2(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G2078), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n786), .C1(new_n754), .C2(new_n760), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT30), .B(G28), .ZN(new_n788));
  OR2_X1    g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  NAND2_X1  g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n788), .A2(new_n719), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n791), .B1(new_n719), .B2(new_n639), .C1(new_n785), .C2(G2078), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n782), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n715), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n752), .A2(new_n753), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n781), .A2(new_n793), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n705), .A2(new_n706), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n762), .A2(new_n763), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n765), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n715), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n715), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT93), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n809), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n715), .A2(G6), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G305), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n715), .A2(G22), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n715), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n814), .B2(new_n813), .ZN(new_n821));
  OR3_X1    g396(.A1(new_n816), .A2(KEYINPUT34), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT34), .B1(new_n816), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n479), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n489), .A2(G119), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n480), .A2(G107), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT90), .Z(new_n829));
  MUX2_X1   g404(.A(G25), .B(new_n829), .S(G29), .Z(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G290), .A2(G16), .ZN(new_n834));
  INV_X1    g409(.A(G24), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n835), .A2(KEYINPUT91), .A3(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT91), .B1(new_n835), .B2(G16), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1986), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n822), .A2(new_n823), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n736), .A2(new_n802), .A3(new_n843), .A4(new_n845), .ZN(G150));
  INV_X1    g421(.A(G150), .ZN(G311));
  AOI22_X1  g422(.A1(new_n536), .A2(G55), .B1(G93), .B2(new_n526), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  INV_X1    g424(.A(G80), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n553), .A2(new_n849), .B1(new_n850), .B2(new_n532), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT104), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n853), .B1(new_n850), .B2(new_n532), .C1(new_n553), .C2(new_n849), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(G651), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n612), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n848), .B2(new_n855), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n848), .A2(new_n855), .A3(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n562), .ZN(new_n866));
  INV_X1    g441(.A(new_n864), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n862), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n563), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n860), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n620), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n858), .B1(new_n873), .B2(new_n874), .ZN(G145));
  XOR2_X1   g450(.A(G160), .B(new_n639), .Z(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n744), .A2(new_n772), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n744), .A2(new_n772), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n479), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n489), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n480), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n828), .B(new_n885), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n879), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n879), .B2(new_n880), .ZN(new_n888));
  XNOR2_X1  g463(.A(G164), .B(new_n726), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(new_n631), .Z(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n878), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n877), .A3(new_n891), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g474(.A1(new_n856), .A2(G868), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n870), .A2(new_n624), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n623), .B1(new_n869), .B2(new_n866), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n611), .A2(G299), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n617), .B1(new_n610), .B2(new_n607), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n612), .A2(new_n617), .ZN(new_n910));
  INV_X1    g485(.A(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT41), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n906), .B2(new_n907), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n902), .A2(new_n904), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(KEYINPUT107), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n905), .A2(new_n908), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n916), .ZN(new_n921));
  XNOR2_X1  g496(.A(G305), .B(G303), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(new_n804), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n925));
  XOR2_X1   g500(.A(new_n924), .B(new_n925), .Z(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n909), .A2(new_n928), .A3(KEYINPUT107), .A4(new_n917), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n900), .B1(new_n930), .B2(G868), .ZN(G295));
  AOI21_X1  g506(.A(new_n900), .B1(new_n930), .B2(G868), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(G301), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(G301), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(G168), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(G171), .A2(KEYINPUT108), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n934), .A3(G286), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n869), .B2(new_n866), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n865), .A2(new_n562), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n868), .A2(new_n563), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n939), .A4(new_n937), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n941), .A2(new_n908), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n912), .A2(new_n914), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n941), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n924), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND4_X1   g523(.A1(new_n943), .A2(new_n942), .A3(new_n939), .A4(new_n937), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n942), .A2(new_n943), .B1(new_n937), .B2(new_n939), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n915), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n924), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n908), .A3(new_n944), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n897), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n924), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n961), .B(new_n962), .ZN(G397));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(G164), .B2(G1384), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n478), .A2(new_n482), .A3(G40), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n726), .B(G2067), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n744), .B2(G1996), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n971), .A2(new_n744), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI221_X1 g551(.A(KEYINPUT110), .B1(new_n969), .B2(new_n973), .C1(new_n971), .C2(new_n744), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n829), .A2(new_n832), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n727), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n969), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT125), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT125), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n985), .B(new_n969), .C1(new_n979), .C2(new_n981), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n971), .B(KEYINPUT46), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n983), .B1(new_n744), .B2(new_n972), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n828), .B(new_n832), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n977), .A3(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT48), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n990), .A2(new_n991), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n984), .A2(new_n986), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1000));
  INV_X1    g575(.A(new_n507), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n506), .B1(new_n628), .B2(new_n503), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n496), .B(new_n500), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1000), .A2(new_n754), .A3(new_n968), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT45), .B(new_n1008), .C1(new_n1009), .C2(new_n501), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n965), .A2(new_n968), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n778), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n967), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n754), .A4(new_n1000), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1007), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT112), .B(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1017), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1018), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1025), .B2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(KEYINPUT121), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1028), .B(new_n1022), .C1(new_n1025), .C2(new_n1023), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1019), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(new_n1019), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1011), .A2(new_n819), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1013), .A2(new_n706), .A3(new_n1000), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT111), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1038), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1020), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1038), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1037), .A2(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G164), .A2(G1384), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1017), .B1(new_n1053), .B2(new_n968), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n804), .B2(G1976), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n804), .A2(G1976), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1054), .B(new_n1055), .C1(KEYINPUT52), .C2(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT114), .B(G1981), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n590), .B(new_n1063), .C1(new_n596), .C2(new_n597), .ZN(new_n1064));
  INV_X1    g639(.A(new_n590), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1065), .B2(new_n594), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1054), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1011), .B2(G2078), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1005), .A2(new_n968), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n753), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1011), .A2(new_n1073), .A3(G2078), .ZN(new_n1080));
  AOI21_X1  g655(.A(G301), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1052), .A2(new_n1072), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1031), .A2(new_n1033), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(KEYINPUT116), .A2(KEYINPUT63), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1062), .B(new_n1071), .C1(new_n1037), .C2(new_n1050), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1016), .A2(G168), .A3(new_n1020), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(KEYINPUT116), .A2(KEYINPUT63), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT49), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1054), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1064), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1088), .B1(new_n1094), .B2(new_n1054), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1047), .A2(new_n1037), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1050), .B1(new_n1048), .B2(new_n1020), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1086), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT63), .B1(new_n1037), .B2(new_n1050), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1072), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1087), .B(new_n1095), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G301), .B(KEYINPUT54), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n967), .A2(KEYINPUT122), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1073), .A2(G2078), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n478), .A2(new_n482), .A3(new_n1106), .A4(G40), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n965), .A2(new_n1010), .ZN(new_n1109));
  OR3_X1    g684(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT123), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1103), .B1(new_n1112), .B2(new_n1079), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1074), .A2(new_n1080), .A3(new_n1103), .A4(new_n1078), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1052), .B(new_n1072), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G299), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n577), .A2(new_n582), .A3(new_n1117), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(G2072), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n965), .A2(new_n1010), .A3(new_n968), .A4(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1121), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1116), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT61), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n967), .A2(G164), .A3(G1384), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(new_n980), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1348), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n612), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n980), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n611), .B(new_n1135), .C1(new_n1136), .C2(G1348), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1138), .A2(KEYINPUT60), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1116), .B(new_n1142), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT58), .B(G1341), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1011), .A2(G1996), .B1(new_n1131), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n563), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n563), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1130), .A2(new_n1141), .A3(new_n1143), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(new_n1128), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1115), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1102), .B1(new_n1155), .B2(new_n1030), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1083), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G290), .B(G1986), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n983), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n976), .A2(new_n977), .A3(new_n1159), .A4(new_n993), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT124), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1163), .B(new_n1160), .C1(new_n1083), .C2(new_n1156), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n999), .B1(new_n1162), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g740(.A1(new_n469), .A2(G227), .ZN(new_n1167));
  NAND4_X1  g741(.A1(new_n898), .A2(new_n659), .A3(new_n701), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n961), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n1171));
  AOI211_X1 g745(.A(new_n1171), .B(new_n1168), .C1(new_n956), .C2(new_n960), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1172), .ZN(G308));
  NOR2_X1   g747(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n1174));
  AOI21_X1  g748(.A(new_n959), .B1(new_n958), .B2(new_n954), .ZN(new_n1175));
  OAI21_X1  g749(.A(new_n1169), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1176), .A2(new_n1171), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n961), .A2(KEYINPUT127), .A3(new_n1169), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1178), .ZN(G225));
endmodule


