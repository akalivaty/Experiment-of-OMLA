

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n532), .ZN(n888) );
  AND2_X2 U552 ( .A1(n524), .A2(G2104), .ZN(n887) );
  NOR2_X1 U553 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U554 ( .A1(n672), .A2(G8), .ZN(n673) );
  INV_X1 U555 ( .A(n937), .ZN(n692) );
  XOR2_X1 U556 ( .A(n605), .B(KEYINPUT99), .Z(n516) );
  NOR2_X1 U557 ( .A1(n693), .A2(n692), .ZN(n517) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n661) );
  XNOR2_X1 U559 ( .A(n662), .B(n661), .ZN(n675) );
  NOR2_X1 U560 ( .A1(G1966), .A2(n705), .ZN(n678) );
  XNOR2_X1 U561 ( .A(n600), .B(KEYINPUT64), .ZN(n624) );
  XNOR2_X1 U562 ( .A(n673), .B(KEYINPUT32), .ZN(n698) );
  INV_X1 U563 ( .A(n602), .ZN(n665) );
  NAND2_X1 U564 ( .A1(n665), .A2(G8), .ZN(n705) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n524), .ZN(n883) );
  NOR2_X1 U567 ( .A1(G651), .A2(n581), .ZN(n782) );
  NOR2_X1 U568 ( .A1(n530), .A2(n529), .ZN(G160) );
  INV_X1 U569 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U570 ( .A1(n883), .A2(G125), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n887), .A2(G101), .ZN(n518) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U573 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT65), .B(n521), .Z(n530) );
  INV_X1 U575 ( .A(KEYINPUT67), .ZN(n528) );
  XOR2_X1 U576 ( .A(KEYINPUT66), .B(n522), .Z(n523) );
  XNOR2_X1 U577 ( .A(KEYINPUT17), .B(n523), .ZN(n531) );
  NAND2_X1 U578 ( .A1(G137), .A2(n531), .ZN(n526) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U580 ( .A1(n884), .A2(G113), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U582 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G102), .A2(n887), .ZN(n534) );
  INV_X1 U584 ( .A(n531), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G138), .A2(n888), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G126), .A2(n883), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G114), .A2(n884), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U590 ( .A1(n538), .A2(n537), .ZN(G164) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n581) );
  NAND2_X1 U592 ( .A1(n782), .A2(G53), .ZN(n542) );
  INV_X1 U593 ( .A(G651), .ZN(n544) );
  NOR2_X1 U594 ( .A1(G543), .A2(n544), .ZN(n539) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n539), .Z(n540) );
  XNOR2_X1 U596 ( .A(KEYINPUT68), .B(n540), .ZN(n787) );
  NAND2_X1 U597 ( .A1(G65), .A2(n787), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U599 ( .A(KEYINPUT73), .B(n543), .ZN(n549) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U601 ( .A1(G91), .A2(n783), .ZN(n546) );
  NOR2_X1 U602 ( .A1(n581), .A2(n544), .ZN(n784) );
  NAND2_X1 U603 ( .A1(G78), .A2(n784), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT72), .B(n547), .Z(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(G299) );
  NAND2_X1 U607 ( .A1(n783), .A2(G90), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT71), .B(n550), .Z(n552) );
  NAND2_X1 U609 ( .A1(n784), .A2(G77), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT9), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G52), .A2(n782), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n787), .A2(G64), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT70), .B(n556), .Z(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n783), .A2(G89), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G76), .A2(n784), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT5), .ZN(n568) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n782), .A2(G51), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G63), .A2(n787), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n566), .B(n565), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(n569), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G88), .A2(n783), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G75), .A2(n784), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n782), .A2(G50), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT88), .B(n572), .Z(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G62), .A2(n787), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(G303) );
  NAND2_X1 U638 ( .A1(G49), .A2(n782), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT86), .B(n579), .ZN(n580) );
  NOR2_X1 U642 ( .A1(n787), .A2(n580), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n581), .A2(G87), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U645 ( .A1(n783), .A2(G86), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G61), .A2(n787), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G73), .A2(n784), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT2), .ZN(n587) );
  XNOR2_X1 U650 ( .A(n587), .B(KEYINPUT87), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n782), .A2(G48), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G85), .A2(n783), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G72), .A2(n784), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G60), .A2(n787), .ZN(n594) );
  XNOR2_X1 U658 ( .A(KEYINPUT69), .B(n594), .ZN(n595) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n782), .A2(G47), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(G290) );
  NAND2_X1 U662 ( .A1(G160), .A2(G40), .ZN(n727) );
  INV_X1 U663 ( .A(n727), .ZN(n599) );
  NOR2_X1 U664 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X1 U665 ( .A1(n599), .A2(n728), .ZN(n600) );
  INV_X1 U666 ( .A(n624), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G2067), .A2(n602), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT98), .ZN(n604) );
  NAND2_X1 U669 ( .A1(G1348), .A2(n665), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U671 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n607) );
  NAND2_X1 U672 ( .A1(G81), .A2(n783), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U674 ( .A1(n784), .A2(G68), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U676 ( .A(KEYINPUT13), .B(n610), .Z(n613) );
  NAND2_X1 U677 ( .A1(n787), .A2(G56), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n611), .Z(n612) );
  NOR2_X1 U679 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U680 ( .A1(n782), .A2(G43), .ZN(n614) );
  NAND2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n921) );
  INV_X1 U682 ( .A(n921), .ZN(n632) );
  NAND2_X1 U683 ( .A1(n783), .A2(G92), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G66), .A2(n787), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G79), .A2(n784), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G54), .A2(n782), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U690 ( .A(KEYINPUT15), .B(n622), .Z(n623) );
  XNOR2_X1 U691 ( .A(KEYINPUT76), .B(n623), .ZN(n800) );
  AND2_X1 U692 ( .A1(n632), .A2(n800), .ZN(n628) );
  INV_X1 U693 ( .A(n624), .ZN(n650) );
  NAND2_X1 U694 ( .A1(n650), .A2(G1996), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT26), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n665), .A2(G1341), .ZN(n626) );
  AND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U698 ( .A1(n628), .A2(n631), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n516), .A2(n629), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT100), .ZN(n635) );
  AND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U702 ( .A1(n800), .A2(n633), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n641) );
  INV_X1 U704 ( .A(G299), .ZN(n643) );
  XOR2_X1 U705 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n637) );
  NAND2_X1 U706 ( .A1(G2072), .A2(n650), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U708 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U709 ( .A1(n650), .A2(n949), .ZN(n638) );
  NOR2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U714 ( .A(n644), .B(KEYINPUT28), .Z(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U716 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n654) );
  NOR2_X1 U718 ( .A1(n650), .A2(G1961), .ZN(n649) );
  XOR2_X1 U719 ( .A(KEYINPUT96), .B(n649), .Z(n652) );
  XNOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .ZN(n1004) );
  NAND2_X1 U721 ( .A1(n650), .A2(n1004), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n658), .A2(G171), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n676) );
  NOR2_X1 U725 ( .A1(n665), .A2(G2084), .ZN(n674) );
  NOR2_X1 U726 ( .A1(n678), .A2(n674), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G8), .A2(n655), .ZN(n656) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n656), .ZN(n657) );
  NOR2_X1 U729 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U730 ( .A1(G171), .A2(n658), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n676), .A2(n675), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n663), .A2(G286), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT102), .ZN(n671) );
  NOR2_X1 U734 ( .A1(n665), .A2(G2090), .ZN(n667) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n705), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n668), .A2(G303), .ZN(n669) );
  XOR2_X1 U738 ( .A(KEYINPUT103), .B(n669), .Z(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U740 ( .A1(G8), .A2(n674), .ZN(n680) );
  AND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n699) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n925) );
  AND2_X1 U745 ( .A1(n699), .A2(n925), .ZN(n681) );
  AND2_X1 U746 ( .A1(n698), .A2(n681), .ZN(n688) );
  INV_X1 U747 ( .A(n925), .ZN(n683) );
  NOR2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NOR2_X1 U749 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n690), .A2(n682), .ZN(n930) );
  OR2_X1 U751 ( .A1(n683), .A2(n930), .ZN(n684) );
  OR2_X1 U752 ( .A1(n705), .A2(n684), .ZN(n686) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  INV_X1 U756 ( .A(n689), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n690), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n691), .A2(n705), .ZN(n693) );
  XOR2_X1 U759 ( .A(G1981), .B(G305), .Z(n937) );
  NAND2_X1 U760 ( .A1(n694), .A2(n517), .ZN(n695) );
  XNOR2_X1 U761 ( .A(n695), .B(KEYINPUT104), .ZN(n709) );
  NOR2_X1 U762 ( .A1(G2090), .A2(G303), .ZN(n696) );
  XOR2_X1 U763 ( .A(KEYINPUT105), .B(n696), .Z(n697) );
  NAND2_X1 U764 ( .A1(G8), .A2(n697), .ZN(n701) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  AND2_X1 U767 ( .A1(n702), .A2(n705), .ZN(n707) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U769 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n744) );
  NAND2_X1 U773 ( .A1(G95), .A2(n887), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G131), .A2(n888), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U776 ( .A(KEYINPUT94), .B(n712), .ZN(n716) );
  NAND2_X1 U777 ( .A1(G119), .A2(n883), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G107), .A2(n884), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n900) );
  INV_X1 U781 ( .A(G1991), .ZN(n997) );
  NOR2_X1 U782 ( .A1(n900), .A2(n997), .ZN(n726) );
  NAND2_X1 U783 ( .A1(G105), .A2(n887), .ZN(n717) );
  XNOR2_X1 U784 ( .A(n717), .B(KEYINPUT38), .ZN(n724) );
  NAND2_X1 U785 ( .A1(G129), .A2(n883), .ZN(n719) );
  NAND2_X1 U786 ( .A1(G117), .A2(n884), .ZN(n718) );
  NAND2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G141), .A2(n888), .ZN(n720) );
  XNOR2_X1 U789 ( .A(KEYINPUT95), .B(n720), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n869) );
  AND2_X1 U792 ( .A1(n869), .A2(G1996), .ZN(n725) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n970) );
  NOR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n753) );
  INV_X1 U795 ( .A(n753), .ZN(n729) );
  NOR2_X1 U796 ( .A1(n970), .A2(n729), .ZN(n747) );
  INV_X1 U797 ( .A(n747), .ZN(n742) );
  XOR2_X1 U798 ( .A(G1986), .B(G290), .Z(n929) );
  NAND2_X1 U799 ( .A1(G128), .A2(n883), .ZN(n731) );
  NAND2_X1 U800 ( .A1(G116), .A2(n884), .ZN(n730) );
  NAND2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U802 ( .A(n732), .B(KEYINPUT35), .ZN(n737) );
  NAND2_X1 U803 ( .A1(G104), .A2(n887), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G140), .A2(n888), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U806 ( .A(KEYINPUT34), .B(n735), .Z(n736) );
  NAND2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U808 ( .A(n738), .B(KEYINPUT36), .Z(n898) );
  XNOR2_X1 U809 ( .A(G2067), .B(KEYINPUT37), .ZN(n751) );
  OR2_X1 U810 ( .A1(n898), .A2(n751), .ZN(n739) );
  XOR2_X1 U811 ( .A(KEYINPUT93), .B(n739), .Z(n977) );
  NAND2_X1 U812 ( .A1(n929), .A2(n977), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n740), .A2(n753), .ZN(n741) );
  AND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n756) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n869), .ZN(n973) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n745) );
  AND2_X1 U818 ( .A1(n997), .A2(n900), .ZN(n988) );
  NOR2_X1 U819 ( .A1(n745), .A2(n988), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n973), .A2(n748), .ZN(n749) );
  XNOR2_X1 U822 ( .A(n749), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n750), .A2(n977), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n751), .A2(n898), .ZN(n987) );
  NAND2_X1 U825 ( .A1(n752), .A2(n987), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U828 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U830 ( .A1(n888), .A2(G135), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n758), .B(KEYINPUT80), .ZN(n766) );
  NAND2_X1 U832 ( .A1(n883), .A2(G123), .ZN(n759) );
  XNOR2_X1 U833 ( .A(n759), .B(KEYINPUT18), .ZN(n761) );
  NAND2_X1 U834 ( .A1(G111), .A2(n884), .ZN(n760) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U836 ( .A1(G99), .A2(n887), .ZN(n762) );
  XNOR2_X1 U837 ( .A(KEYINPUT81), .B(n762), .ZN(n763) );
  NOR2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n986) );
  XNOR2_X1 U840 ( .A(G2096), .B(n986), .ZN(n767) );
  OR2_X1 U841 ( .A1(G2100), .A2(n767), .ZN(G156) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n822) );
  NAND2_X1 U847 ( .A1(n822), .A2(G567), .ZN(n769) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n774) );
  OR2_X1 U850 ( .A1(n921), .A2(n774), .ZN(G153) );
  INV_X1 U851 ( .A(G171), .ZN(G301) );
  INV_X1 U852 ( .A(G868), .ZN(n804) );
  NOR2_X1 U853 ( .A1(G301), .A2(n804), .ZN(n771) );
  INV_X1 U854 ( .A(n800), .ZN(n926) );
  NOR2_X1 U855 ( .A1(n926), .A2(G868), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(G284) );
  NOR2_X1 U857 ( .A1(G286), .A2(n804), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n775), .A2(n800), .ZN(n776) );
  XNOR2_X1 U862 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U863 ( .A1(G868), .A2(n800), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G559), .A2(n777), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT78), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n921), .A2(G868), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U868 ( .A(KEYINPUT79), .B(n781), .Z(G282) );
  INV_X1 U869 ( .A(G303), .ZN(G166) );
  NAND2_X1 U870 ( .A1(G55), .A2(n782), .ZN(n792) );
  NAND2_X1 U871 ( .A1(G93), .A2(n783), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n787), .A2(G67), .ZN(n788) );
  XOR2_X1 U875 ( .A(KEYINPUT84), .B(n788), .Z(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U878 ( .A(n793), .B(KEYINPUT85), .ZN(n919) );
  XNOR2_X1 U879 ( .A(n919), .B(G299), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n794), .B(G288), .ZN(n795) );
  XOR2_X1 U881 ( .A(n795), .B(KEYINPUT19), .Z(n797) );
  XNOR2_X1 U882 ( .A(G166), .B(KEYINPUT89), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n798), .B(G305), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(G290), .ZN(n904) );
  XNOR2_X1 U886 ( .A(n921), .B(KEYINPUT82), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n800), .A2(G559), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n802), .B(n801), .ZN(n916) );
  XNOR2_X1 U889 ( .A(n904), .B(n916), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n803), .A2(G868), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n804), .A2(n919), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U893 ( .A(KEYINPUT90), .B(n807), .Z(G295) );
  NAND2_X1 U894 ( .A1(G2078), .A2(G2084), .ZN(n808) );
  XOR2_X1 U895 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U896 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U897 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XOR2_X1 U899 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U901 ( .A1(G120), .A2(G69), .ZN(n812) );
  NOR2_X1 U902 ( .A1(G237), .A2(n812), .ZN(n813) );
  XNOR2_X1 U903 ( .A(KEYINPUT92), .B(n813), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(G108), .ZN(n914) );
  NAND2_X1 U905 ( .A1(n914), .A2(G567), .ZN(n820) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n816) );
  XNOR2_X1 U907 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n815) );
  XNOR2_X1 U908 ( .A(n816), .B(n815), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n817), .A2(G218), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G96), .A2(n818), .ZN(n915) );
  NAND2_X1 U911 ( .A1(n915), .A2(G2106), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n920) );
  NAND2_X1 U913 ( .A1(G483), .A2(G661), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n920), .A2(n821), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n822), .ZN(G217) );
  INV_X1 U917 ( .A(G661), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G2), .A2(G15), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U920 ( .A(KEYINPUT108), .B(n825), .Z(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G2454), .B(G2435), .ZN(n836) );
  XNOR2_X1 U924 ( .A(KEYINPUT106), .B(G2427), .ZN(n834) );
  XOR2_X1 U925 ( .A(G2430), .B(G2446), .Z(n829) );
  XNOR2_X1 U926 ( .A(G2443), .B(G2451), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n830), .B(G2438), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1341), .B(G1348), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n837), .A2(G14), .ZN(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT107), .B(n838), .ZN(G401) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2090), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2072), .B(G2084), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U938 ( .A(n841), .B(G2100), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2078), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n845) );
  XNOR2_X1 U942 ( .A(KEYINPUT109), .B(G2678), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U945 ( .A(G1991), .B(G1976), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1971), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n859) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G2474), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1956), .B(KEYINPUT110), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(G1986), .B(G1981), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G100), .A2(n887), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n860), .B(KEYINPUT114), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n862) );
  NAND2_X1 U961 ( .A1(G124), .A2(n883), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n884), .A2(G112), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G136), .A2(n888), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(G162) );
  XNOR2_X1 U968 ( .A(G162), .B(n869), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n870), .B(n986), .ZN(n874) );
  XOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n872) );
  XNOR2_X1 U971 ( .A(G164), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U973 ( .A(n874), .B(n873), .Z(n897) );
  NAND2_X1 U974 ( .A1(G103), .A2(n887), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G139), .A2(n888), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G127), .A2(n883), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G115), .A2(n884), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT116), .B(n882), .Z(n979) );
  NAND2_X1 U983 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G106), .A2(n887), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G142), .A2(n888), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(KEYINPUT115), .B(n891), .ZN(n892) );
  XNOR2_X1 U990 ( .A(KEYINPUT45), .B(n892), .ZN(n893) );
  NOR2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n979), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n902) );
  XNOR2_X1 U995 ( .A(G160), .B(n900), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U998 ( .A(n904), .B(G286), .Z(n906) );
  XNOR2_X1 U999 ( .A(n926), .B(G171), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n907), .B(n921), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G397) );
  OR2_X1 U1003 ( .A1(n920), .A2(G401), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G225) );
  XOR2_X1 U1009 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  NOR2_X1 U1017 ( .A1(n916), .A2(G860), .ZN(n917) );
  XOR2_X1 U1018 ( .A(KEYINPUT83), .B(n917), .Z(n918) );
  XNOR2_X1 U1019 ( .A(n919), .B(n918), .ZN(G145) );
  INV_X1 U1020 ( .A(n920), .ZN(G319) );
  XNOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .ZN(n943) );
  XOR2_X1 U1022 ( .A(n921), .B(G1341), .Z(n923) );
  XNOR2_X1 U1023 ( .A(G171), .B(G1961), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n936) );
  NAND2_X1 U1025 ( .A1(G1971), .A2(G303), .ZN(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G1348), .B(n926), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(G1966), .B(G168), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(KEYINPUT57), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n1025) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT125), .ZN(n968) );
  XNOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(G4), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n952) );
  XOR2_X1 U1046 ( .A(KEYINPUT126), .B(n949), .Z(n950) );
  XNOR2_X1 U1047 ( .A(G20), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n953), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n961) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1061 ( .A(n965), .B(KEYINPUT61), .Z(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT127), .B(n966), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n969), .A2(G11), .ZN(n1023) );
  INV_X1 U1065 ( .A(G29), .ZN(n1019) );
  XNOR2_X1 U1066 ( .A(G160), .B(G2084), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n976) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT51), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n985) );
  XOR2_X1 U1073 ( .A(G2072), .B(n979), .Z(n981) );
  XNOR2_X1 U1074 ( .A(G2078), .B(G164), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT50), .B(n982), .Z(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(n983), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT52), .B(n992), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT120), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(KEYINPUT55), .A2(n994), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n1019), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT121), .ZN(n1021) );
  XOR2_X1 U1087 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n1017) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G35), .ZN(n1012) );
  XNOR2_X1 U1089 ( .A(G25), .B(n997), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(G2067), .B(G26), .Z(n998) );
  NAND2_X1 U1091 ( .A1(n998), .A2(G28), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G33), .B(G2072), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n999), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(n1004), .B(G27), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(G1996), .B(G32), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1099 ( .A(n1007), .B(KEYINPUT123), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(KEYINPUT53), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(G2084), .B(G34), .Z(n1013) );
  XNOR2_X1 U1104 ( .A(KEYINPUT54), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

