//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G125), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT69), .A4(G125), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n194), .A2(new_n198), .A3(G146), .A4(new_n199), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT70), .A3(new_n201), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(G237), .A2(G953), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT85), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT85), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(G214), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G214), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT85), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n211), .B2(new_n214), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(KEYINPUT17), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n207), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n195), .A2(new_n197), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n201), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n195), .A2(new_n197), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n217), .A2(KEYINPUT18), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n211), .B(new_n214), .C1(new_n226), .C2(new_n215), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n227), .A2(KEYINPUT86), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(KEYINPUT86), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT87), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n208), .A2(G214), .B1(KEYINPUT85), .B2(G143), .ZN(new_n232));
  INV_X1    g046(.A(new_n212), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT85), .B(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n235), .B(new_n236), .C1(new_n226), .C2(new_n215), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n227), .A2(KEYINPUT86), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT87), .B1(new_n239), .B2(new_n225), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n189), .B(new_n220), .C1(new_n231), .C2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n204), .B1(new_n216), .B2(new_n217), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n243));
  XOR2_X1   g057(.A(new_n243), .B(KEYINPUT19), .Z(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n244), .B2(new_n201), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n248), .B2(new_n230), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n241), .B1(new_n249), .B2(new_n189), .ZN(new_n250));
  NOR2_X1   g064(.A1(G475), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT20), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n243), .B(KEYINPUT19), .ZN(new_n255));
  OAI221_X1 g069(.A(new_n204), .B1(new_n216), .B2(new_n217), .C1(new_n255), .C2(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n231), .B2(new_n240), .ZN(new_n257));
  INV_X1    g071(.A(new_n189), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n254), .B1(new_n259), .B2(new_n241), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G478), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT15), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT9), .B(G234), .ZN(new_n267));
  INV_X1    g081(.A(G217), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n267), .A2(new_n268), .A3(G953), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G116), .B(G122), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(G107), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT89), .ZN(new_n273));
  XOR2_X1   g087(.A(G116), .B(G122), .Z(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G107), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT89), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT13), .B1(new_n281), .B2(G143), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G128), .B(G143), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n273), .A2(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n290));
  OAI211_X1 g104(.A(G107), .B(new_n290), .C1(new_n274), .C2(KEYINPUT14), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(G134), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n285), .A2(G134), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n291), .A2(new_n277), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n270), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n287), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n272), .A2(KEYINPUT89), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n278), .A2(new_n279), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n294), .A3(new_n269), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n266), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(G902), .B(new_n265), .C1(new_n296), .C2(new_n301), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G953), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n307), .A2(G952), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT90), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n220), .B1(new_n231), .B2(new_n240), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n258), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n241), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n303), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G475), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n263), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G143), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT1), .B1(new_n323), .B2(G146), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(G146), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n201), .A2(G143), .ZN(new_n326));
  OAI211_X1 g140(.A(G128), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n201), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(G146), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(new_n329), .C1(KEYINPUT1), .C2(new_n281), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n196), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n333));
  XNOR2_X1  g147(.A(G143), .B(G146), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT0), .B(G128), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT0), .A2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n329), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT0), .A2(G128), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT64), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n332), .B1(new_n343), .B2(new_n196), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT82), .B(G224), .Z(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT7), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n350));
  INV_X1    g164(.A(G119), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G116), .ZN(new_n352));
  XNOR2_X1  g166(.A(G116), .B(G119), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(G113), .B(new_n352), .C1(new_n354), .C2(new_n350), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT2), .B(G113), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n353), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n188), .B2(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n276), .A2(KEYINPUT3), .A3(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT77), .B1(new_n276), .B2(G104), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n188), .A3(G107), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n276), .B2(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n276), .A2(G104), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n188), .A2(KEYINPUT78), .A3(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G101), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n355), .A2(new_n358), .A3(new_n367), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G122), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n276), .A2(KEYINPUT3), .A3(G104), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n276), .B2(G104), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n364), .A2(new_n366), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n354), .A2(new_n356), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n358), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(G101), .C1(new_n378), .C2(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n375), .C1(new_n381), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n355), .A2(new_n358), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n367), .A2(new_n373), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n374), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n375), .B(KEYINPUT8), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n344), .A2(new_n348), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n349), .A2(new_n387), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n303), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n374), .B1(new_n381), .B2(new_n386), .ZN(new_n397));
  INV_X1    g211(.A(new_n375), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n387), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n383), .A3(new_n385), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n375), .B1(new_n403), .B2(new_n374), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n406), .A3(new_n398), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n400), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n344), .B(new_n347), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n396), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n413), .B(new_n414), .C1(KEYINPUT83), .C2(new_n416), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n410), .A2(new_n412), .ZN(new_n420));
  INV_X1    g234(.A(new_n396), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT84), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n267), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n307), .A2(G227), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n283), .B2(G137), .ZN(new_n434));
  INV_X1    g248(.A(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT11), .A3(G134), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n283), .A2(G137), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n436), .A3(new_n215), .A4(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n402), .A2(new_n343), .A3(new_n385), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n367), .A2(new_n373), .A3(new_n330), .A4(new_n327), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT10), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n327), .A2(new_n330), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(KEYINPUT10), .A3(new_n367), .A4(new_n373), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n441), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n402), .A2(new_n343), .A3(new_n385), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n445), .A3(new_n447), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n441), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n439), .A2(new_n440), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n451), .A2(new_n456), .A3(new_n445), .A4(new_n447), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n432), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n389), .A2(new_n331), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n443), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT79), .A3(new_n441), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT12), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n460), .A2(KEYINPUT79), .A3(new_n463), .A4(new_n441), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n457), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n465), .A2(new_n466), .A3(new_n431), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n428), .B(new_n303), .C1(new_n458), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n428), .A2(new_n303), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n466), .A2(new_n431), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n457), .A3(new_n464), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n455), .A2(new_n470), .B1(new_n431), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n472), .B2(G469), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n427), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n322), .A2(new_n424), .A3(new_n425), .A4(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT32), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT31), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n383), .B(KEYINPUT66), .ZN(new_n479));
  INV_X1    g293(.A(new_n437), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n283), .A2(G137), .ZN(new_n481));
  OAI21_X1  g295(.A(G131), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(new_n327), .A3(new_n440), .A4(new_n330), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n456), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(KEYINPUT65), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(KEYINPUT65), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n441), .A2(new_n336), .A3(new_n338), .A4(new_n342), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n491), .A2(KEYINPUT65), .A3(new_n487), .A4(new_n483), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n493), .B2(new_n383), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n208), .A2(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n478), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n383), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n490), .B2(new_n492), .ZN(new_n501));
  INV_X1    g315(.A(new_n498), .ZN(new_n502));
  NOR4_X1   g316(.A1(new_n501), .A2(KEYINPUT31), .A3(new_n486), .A4(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT28), .B1(new_n479), .B2(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(new_n485), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n383), .B(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n485), .A2(new_n383), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n498), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n499), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n477), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n512), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n493), .A2(new_n383), .ZN(new_n518));
  INV_X1    g332(.A(new_n486), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n498), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT31), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n494), .A2(new_n478), .A3(new_n498), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT32), .A3(new_n514), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n505), .A2(new_n508), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n504), .B2(new_n509), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n502), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n510), .A2(new_n511), .A3(new_n498), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n527), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n494), .A2(new_n498), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n516), .A2(new_n524), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G110), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT24), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G110), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G119), .B(G128), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n545));
  OAI211_X1 g359(.A(G119), .B(new_n281), .C1(new_n545), .C2(KEYINPUT23), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n351), .B2(G128), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT68), .B1(new_n351), .B2(G128), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n543), .A2(new_n544), .B1(G110), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n205), .A2(new_n206), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n543), .A2(new_n544), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT71), .B(G110), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n204), .B(new_n222), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT72), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT22), .B(G137), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n552), .A2(new_n556), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n268), .B1(G234), .B2(new_n303), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT75), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT73), .B1(new_n570), .B2(KEYINPUT25), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n552), .A2(new_n556), .A3(new_n561), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n561), .B1(new_n552), .B2(new_n556), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n303), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT74), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n577), .A3(KEYINPUT25), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n579), .A3(new_n575), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n571), .A2(new_n576), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n569), .B1(new_n566), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n476), .B1(new_n535), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n535), .A2(new_n582), .A3(new_n476), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n475), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n363), .ZN(G3));
  NAND2_X1  g401(.A1(new_n523), .A2(new_n303), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT91), .A3(G472), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT91), .A2(G472), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n523), .A2(new_n303), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n474), .A3(new_n582), .A4(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n425), .ZN(new_n594));
  INV_X1    g408(.A(new_n416), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n408), .B(new_n407), .C1(new_n401), .C2(new_n404), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n411), .B1(new_n596), .B2(new_n400), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n597), .B2(new_n396), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n422), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n314), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n264), .A2(new_n303), .ZN(new_n602));
  INV_X1    g416(.A(new_n302), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(new_n264), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n302), .A2(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n302), .A2(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(G478), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI211_X1 g424(.A(KEYINPUT20), .B(new_n254), .C1(new_n259), .C2(new_n241), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n261), .B1(new_n250), .B2(new_n251), .ZN(new_n612));
  INV_X1    g426(.A(G475), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n317), .B2(new_n241), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n601), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n593), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  NAND2_X1  g434(.A1(new_n320), .A2(new_n306), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n612), .B1(new_n611), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n260), .B2(new_n261), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n601), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n593), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  AND3_X1   g445(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n594), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n588), .B(new_n590), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n557), .B1(KEYINPUT36), .B2(new_n561), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n561), .A2(KEYINPUT36), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n552), .A3(new_n556), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n567), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT93), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n581), .B2(new_n566), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n321), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n633), .A2(new_n474), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AND2_X1   g459(.A1(new_n535), .A2(new_n474), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n304), .A2(new_n305), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n319), .B2(G475), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n311), .B(KEYINPUT94), .Z(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n313), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n250), .A2(new_n622), .A3(new_n261), .A4(new_n251), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n253), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n648), .B(new_n653), .C1(new_n655), .C2(new_n624), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n597), .A2(new_n396), .A3(new_n595), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n425), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n656), .A2(new_n659), .A3(new_n641), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n646), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XNOR2_X1  g476(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n424), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n519), .A2(new_n502), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n303), .B1(new_n666), .B2(new_n525), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n494), .A2(new_n502), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n516), .A2(new_n524), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT96), .Z(new_n671));
  XOR2_X1   g485(.A(new_n652), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n474), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n647), .B1(new_n263), .B2(new_n320), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n425), .A3(new_n641), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n665), .A2(new_n671), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  AOI21_X1  g494(.A(new_n609), .B1(new_n263), .B2(new_n320), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n581), .A2(new_n566), .ZN(new_n682));
  INV_X1    g496(.A(new_n640), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n684), .A3(new_n599), .A4(new_n653), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n535), .A2(new_n474), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT97), .B(G146), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G48));
  OAI21_X1  g503(.A(new_n303), .B1(new_n458), .B2(new_n467), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n426), .A3(new_n468), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n535), .A3(new_n582), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n617), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n628), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  NAND4_X1  g512(.A1(new_n599), .A2(new_n426), .A3(new_n468), .A4(new_n691), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n535), .A3(new_n642), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  OAI211_X1 g516(.A(new_n521), .B(new_n522), .C1(new_n498), .C2(new_n526), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n514), .B(KEYINPUT98), .Z(new_n704));
  AOI22_X1  g518(.A1(new_n588), .A2(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n582), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n422), .A2(new_n598), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n615), .A3(new_n425), .A4(new_n306), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n600), .A3(new_n692), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT99), .B(G122), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n681), .A3(new_n684), .A4(new_n653), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n699), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n196), .ZN(G27));
  NAND4_X1  g529(.A1(new_n632), .A2(KEYINPUT100), .A3(new_n425), .A4(new_n474), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n418), .A2(new_n423), .A3(new_n419), .A4(new_n425), .ZN(new_n718));
  INV_X1    g532(.A(new_n474), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n535), .A2(new_n582), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n722), .B1(new_n535), .B2(new_n582), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n610), .A2(new_n615), .A3(new_n653), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n535), .A2(new_n582), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n716), .B2(new_n720), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(KEYINPUT42), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n728), .A2(KEYINPUT42), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  INV_X1    g547(.A(new_n729), .ZN(new_n734));
  INV_X1    g548(.A(new_n656), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n721), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n455), .A2(new_n470), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n471), .A2(new_n431), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n428), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n472), .A2(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n469), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n753), .A3(KEYINPUT46), .A4(new_n747), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n752), .A3(new_n468), .A4(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(new_n426), .A3(new_n672), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n615), .B2(new_n609), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT43), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n634), .A2(new_n641), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n759), .B2(new_n760), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n718), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NOR4_X1   g581(.A1(new_n718), .A2(new_n535), .A3(new_n726), .A4(new_n582), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n426), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT47), .B1(new_n755), .B2(new_n426), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NAND2_X1  g586(.A1(new_n759), .A2(new_n649), .ZN(new_n773));
  INV_X1    g587(.A(new_n718), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n692), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n725), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n582), .A2(new_n311), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n671), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(new_n616), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n759), .A2(new_n649), .A3(new_n706), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n700), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n308), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n769), .A2(new_n770), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n691), .A2(new_n468), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n426), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n774), .B(new_n784), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n692), .A2(new_n594), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n664), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT114), .B1(new_n793), .B2(new_n783), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n784), .A2(new_n796), .A3(new_n664), .A4(new_n792), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n784), .A2(KEYINPUT50), .A3(new_n664), .A4(new_n792), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(KEYINPUT115), .A3(new_n795), .A4(new_n797), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n588), .A2(G472), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n703), .A2(new_n704), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n684), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n773), .A2(new_n806), .A3(new_n775), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT116), .Z(new_n808));
  OR3_X1    g622(.A1(new_n781), .A2(new_n615), .A3(new_n610), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n790), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n786), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT106), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n634), .A2(new_n425), .A3(new_n424), .A4(new_n474), .ZN(new_n815));
  INV_X1    g629(.A(new_n642), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n263), .A2(new_n320), .A3(new_n306), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n616), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n425), .A3(new_n424), .A4(new_n600), .ZN(new_n819));
  OAI22_X1  g633(.A1(new_n815), .A2(new_n816), .B1(new_n819), .B2(new_n592), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n814), .B1(new_n820), .B2(new_n586), .ZN(new_n821));
  INV_X1    g635(.A(new_n475), .ZN(new_n822));
  INV_X1    g636(.A(new_n585), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n823), .B2(new_n583), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n593), .A2(new_n633), .A3(new_n600), .A4(new_n818), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(KEYINPUT106), .A3(new_n825), .A4(new_n643), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n806), .A2(new_n726), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n721), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n306), .A2(new_n652), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n320), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n641), .B(new_n831), .C1(new_n625), .C2(new_n623), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n646), .A3(new_n774), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n736), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n694), .A2(new_n697), .A3(new_n701), .A4(new_n710), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n827), .A2(new_n834), .A3(new_n732), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n700), .A2(new_n828), .B1(new_n646), .B2(new_n660), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n726), .A2(new_n659), .A3(new_n641), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n468), .A2(new_n473), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n653), .A2(KEYINPUT107), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n653), .A2(KEYINPUT107), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n426), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n641), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n708), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n646), .A2(new_n839), .B1(new_n846), .B2(new_n670), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n838), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n626), .A2(new_n599), .A3(new_n684), .A4(new_n653), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n851), .A2(new_n686), .B1(new_n713), .B2(new_n699), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n843), .B1(new_n468), .B2(new_n473), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n675), .A2(new_n853), .A3(new_n599), .A4(new_n641), .ZN(new_n854));
  INV_X1    g668(.A(new_n670), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n686), .A2(new_n685), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n849), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n850), .B1(new_n849), .B2(new_n857), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT110), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n848), .B1(new_n838), .B2(new_n847), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n852), .A2(new_n856), .A3(KEYINPUT109), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT52), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n849), .A2(new_n857), .A3(new_n850), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n837), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n834), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n838), .A2(new_n847), .A3(KEYINPUT52), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT108), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n838), .A2(new_n847), .A3(KEYINPUT108), .A4(KEYINPUT52), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n730), .A2(new_n731), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n835), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n732), .A2(KEYINPUT111), .A3(new_n835), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n872), .A2(new_n877), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT110), .B1(new_n858), .B2(new_n859), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n864), .A2(new_n861), .A3(new_n865), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n836), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n871), .B(new_n884), .C1(new_n888), .C2(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT112), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n837), .A2(new_n868), .A3(new_n877), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(KEYINPUT54), .C1(new_n888), .C2(new_n868), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n885), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n813), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n582), .A2(new_n425), .A3(new_n426), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n615), .A3(new_n609), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n896), .A2(new_n664), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n671), .B2(new_n900), .ZN(G75));
  OAI21_X1  g715(.A(new_n884), .B1(new_n888), .B2(KEYINPUT53), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(G210), .A3(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n410), .B(KEYINPUT118), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n411), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n307), .A2(G952), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n903), .B2(KEYINPUT119), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(KEYINPUT119), .B2(new_n903), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n908), .B(new_n909), .C1(new_n911), .C2(new_n906), .ZN(G51));
  NAND2_X1  g726(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n889), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n469), .B(KEYINPUT57), .Z(new_n916));
  OAI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(new_n458), .B2(new_n467), .ZN(new_n917));
  INV_X1    g731(.A(new_n902), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n918), .A2(new_n303), .A3(new_n746), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n909), .B1(new_n917), .B2(new_n919), .ZN(G54));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n303), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n259), .A3(new_n241), .ZN(new_n923));
  INV_X1    g737(.A(new_n909), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .A4(new_n250), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G60));
  XNOR2_X1  g740(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(new_n602), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n890), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n892), .B1(new_n889), .B2(KEYINPUT112), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n606), .A2(new_n607), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n928), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n909), .B1(new_n914), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n893), .B2(new_n929), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n871), .B1(new_n869), .B2(new_n884), .ZN(new_n941));
  INV_X1    g755(.A(new_n889), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n924), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT121), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n939), .A2(new_n945), .ZN(G63));
  AND2_X1   g760(.A1(new_n635), .A2(new_n637), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n902), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n924), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT61), .B1(new_n952), .B2(KEYINPUT122), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n918), .A2(new_n949), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n924), .B(new_n951), .C1(new_n954), .C2(new_n565), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G66));
  NAND2_X1  g770(.A1(new_n827), .A2(new_n835), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n307), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT123), .Z(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n345), .B2(new_n312), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n904), .B1(G898), .B2(new_n307), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NOR2_X1   g777(.A1(new_n852), .A2(new_n687), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n679), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n774), .A2(new_n474), .A3(new_n672), .A4(new_n818), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n584), .B2(new_n585), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n756), .B2(new_n765), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n771), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n307), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n493), .B(new_n255), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n307), .B1(G227), .B2(G900), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n723), .A2(new_n724), .A3(new_n708), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n756), .B1(new_n765), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n732), .A2(new_n736), .A3(new_n964), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n771), .A2(new_n977), .A3(new_n978), .A4(new_n307), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n974), .A2(KEYINPUT124), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT124), .B1(new_n974), .B2(new_n981), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n979), .A2(new_n980), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n974), .A2(new_n984), .A3(KEYINPUT125), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n975), .B1(new_n984), .B2(KEYINPUT125), .ZN(new_n986));
  OAI22_X1  g800(.A1(new_n982), .A2(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  OAI221_X1 g803(.A(new_n989), .B1(new_n985), .B2(new_n986), .C1(new_n983), .C2(new_n982), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(G72));
  OR2_X1    g805(.A1(new_n971), .A2(new_n957), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  AOI211_X1 g808(.A(new_n502), .B(new_n494), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n771), .A2(new_n977), .A3(new_n978), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n994), .B1(new_n997), .B2(new_n957), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n666), .A2(new_n501), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n909), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n891), .B1(new_n888), .B2(new_n868), .ZN(new_n1001));
  INV_X1    g815(.A(new_n520), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n994), .B1(new_n1002), .B2(new_n532), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n996), .A2(new_n1004), .ZN(G57));
endmodule


