//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n463), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n474), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n474), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n467), .A2(G138), .A3(new_n468), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n462), .A2(new_n464), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n474), .B2(new_n497), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(KEYINPUT69), .B(KEYINPUT4), .C1(new_n474), .C2(new_n497), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(G164));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(new_n508), .A2(new_n512), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G89), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n512), .A2(G543), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT70), .B(G51), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n508), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n510), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n513), .A2(new_n537), .B1(new_n515), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n510), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n513), .A2(new_n543), .B1(new_n515), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  AOI22_X1  g126(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n510), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n513), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n522), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  AND2_X1   g138(.A1(new_n532), .A2(new_n533), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n558), .A2(G87), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n508), .A2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n522), .B2(G49), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G288));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n506), .B2(new_n507), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n575), .B1(new_n571), .B2(new_n572), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n522), .A2(G48), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n555), .A2(G86), .A3(new_n557), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n510), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n513), .A2(new_n584), .B1(new_n515), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n510), .B1(new_n594), .B2(new_n515), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n558), .A2(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n558), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G286), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(G299), .B(KEYINPUT77), .Z(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G297));
  AOI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G280));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n599), .ZN(new_n608));
  INV_X1    g183(.A(new_n595), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G860), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(G559), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT78), .Z(G148));
  OAI21_X1  g188(.A(new_n603), .B1(new_n542), .B2(new_n545), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n610), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n465), .A2(new_n477), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n481), .A2(G123), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT79), .Z(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(new_n469), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n483), .B2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n621), .A2(new_n630), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(KEYINPUT82), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n645), .A2(new_n651), .A3(new_n648), .A4(new_n646), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n647), .B2(new_n649), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT83), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n677), .A3(new_n675), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n680), .A2(new_n682), .A3(new_n683), .A4(new_n685), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n687), .B2(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n671), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n670), .A3(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G23), .B(G288), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT86), .B(G16), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT88), .Z(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AND4_X1   g288(.A1(new_n702), .A2(new_n705), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NOR2_X1   g292(.A1(G25), .A2(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G131), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT85), .Z(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G107), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n625), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n481), .B2(G119), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n707), .A2(G24), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n590), .B2(new_n707), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1986), .Z(new_n731));
  NAND4_X1  g306(.A1(new_n716), .A2(new_n717), .A3(new_n728), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT95), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT94), .B(KEYINPUT25), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n483), .A2(G139), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  AOI22_X1  g314(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(new_n469), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n737), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n743), .B2(G33), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n481), .A2(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n483), .A2(G140), .ZN(new_n752));
  OAI221_X1 g327(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT93), .B(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n706), .A2(G20), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT23), .Z(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G299), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1956), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n745), .A2(new_n746), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n747), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G162), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G35), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT29), .B(G2090), .Z(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT99), .B(G2078), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n771), .B(new_n772), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n707), .A2(G19), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n546), .B2(new_n707), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT90), .B(G1341), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G5), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G301), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n743), .B1(new_n788), .B2(G28), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n790), .A2(KEYINPUT98), .B1(new_n788), .B2(G28), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n785), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n629), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n780), .B(new_n794), .C1(G29), .C2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G4), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n610), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT89), .B(G1348), .Z(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G21), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G168), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1966), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n796), .A2(new_n801), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n743), .A2(G32), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n481), .A2(G129), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT26), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n812), .A2(new_n813), .B1(G105), .B2(new_n477), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n483), .A2(G141), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n808), .B1(new_n817), .B2(new_n743), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT24), .B(G34), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(new_n743), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT97), .Z(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n479), .B2(new_n743), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G2084), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n774), .A2(new_n775), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n820), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n767), .A2(new_n776), .A3(new_n807), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n733), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  AOI22_X1  g405(.A1(G93), .A2(new_n519), .B1(new_n522), .B2(G55), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n510), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n600), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n833), .B(new_n546), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT100), .Z(new_n844));
  OAI21_X1  g419(.A(new_n611), .B1(new_n842), .B2(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n836), .B1(new_n844), .B2(new_n845), .ZN(G145));
  INV_X1    g421(.A(new_n619), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n725), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n483), .A2(G142), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT103), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n481), .A2(G130), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT104), .ZN(new_n852));
  OAI221_X1 g427(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n847), .B1(new_n720), .B2(new_n724), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n848), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n720), .A2(new_n724), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n619), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n854), .B1(new_n860), .B2(new_n856), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n758), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G164), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n501), .A2(new_n502), .ZN(new_n868));
  INV_X1    g443(.A(new_n500), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n504), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n496), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n758), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n742), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n817), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n867), .A2(new_n742), .A3(new_n873), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n865), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(G162), .A2(G160), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n490), .A2(new_n479), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n883), .A3(new_n885), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n795), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n795), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n876), .A2(new_n878), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n817), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n864), .A3(new_n879), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n882), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n891), .B1(new_n882), .B2(new_n894), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(G395));
  INV_X1    g476(.A(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n610), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n600), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n600), .A2(KEYINPUT107), .A3(G299), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT107), .B1(new_n600), .B2(G299), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT108), .B1(new_n905), .B2(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n615), .B(new_n840), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n916), .A2(new_n906), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(G305), .ZN(new_n924));
  XNOR2_X1  g499(.A(G288), .B(G303), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n921), .A2(new_n922), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n833), .A2(new_n603), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n933), .ZN(G331));
  NAND2_X1  g510(.A1(G168), .A2(G171), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G168), .A2(G171), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n840), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n839), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n908), .A2(new_n913), .A3(new_n914), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n906), .A2(new_n941), .A3(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n930), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n928), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n896), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n928), .B1(new_n943), .B2(new_n944), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n911), .A2(new_n942), .A3(KEYINPUT41), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n928), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n905), .B1(new_n942), .B2(KEYINPUT41), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n896), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n951), .A2(new_n955), .A3(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n951), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(KEYINPUT44), .B2(new_n959), .ZN(G397));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G164), .B2(G1384), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n470), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT112), .Z(new_n967));
  XNOR2_X1  g542(.A(new_n758), .B(G2067), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n877), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n966), .A2(G1996), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT46), .Z(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n817), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT111), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n817), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n968), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n975), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n725), .A2(new_n727), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n725), .A2(new_n727), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n967), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n981), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G2067), .B2(new_n758), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n967), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT55), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n872), .A2(KEYINPUT115), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G164), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n872), .A2(new_n993), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n964), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(G2090), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n962), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(KEYINPUT113), .A3(new_n961), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n1007), .B2(new_n965), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1002), .B1(new_n1008), .B2(KEYINPUT114), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n964), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1010), .A2(new_n1011), .A3(G1971), .ZN(new_n1012));
  OAI211_X1 g587(.A(G8), .B(new_n992), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n997), .B1(new_n994), .B2(new_n996), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n965), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(G2090), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n991), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n994), .A2(new_n996), .A3(new_n965), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(G8), .C1(new_n1020), .C2(G288), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G288), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(G1976), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1019), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT116), .B(G1981), .Z(new_n1029));
  NAND4_X1  g604(.A1(new_n580), .A2(new_n577), .A3(new_n578), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT117), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT118), .B(G86), .Z(new_n1032));
  OAI21_X1  g607(.A(new_n579), .B1(new_n513), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G1981), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1028), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1025), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n994), .B2(new_n996), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1003), .A2(new_n965), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n804), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2084), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n998), .A2(new_n1000), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G286), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1013), .A2(new_n1018), .A3(new_n1041), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n991), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1048), .A2(new_n1051), .A3(G286), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1013), .A3(new_n1041), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1013), .A2(new_n1018), .A3(new_n1041), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1043), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2078), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n994), .A2(new_n996), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1059), .B(new_n1061), .C1(new_n1062), .C2(KEYINPUT45), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n998), .A2(new_n1000), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n784), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT124), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1007), .A2(new_n965), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(G2078), .ZN(new_n1073));
  AOI21_X1  g648(.A(G301), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  OAI22_X1  g650(.A1(G168), .A2(new_n1027), .B1(KEYINPUT123), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(KEYINPUT123), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1048), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1078), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1027), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1076), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1047), .A2(G8), .A3(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT62), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1079), .A2(new_n1082), .A3(new_n1086), .A4(new_n1083), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1058), .A2(new_n1074), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1013), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1039), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1031), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1089), .A2(new_n1041), .B1(new_n1028), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1057), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1010), .A2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(G299), .B(KEYINPUT57), .Z(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT119), .B(G1956), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G2067), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n800), .A2(new_n1064), .B1(new_n1026), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n610), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n610), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n610), .B1(new_n1102), .B2(KEYINPUT60), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1106), .A2(new_n1107), .B1(KEYINPUT60), .B2(new_n1102), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT61), .B1(new_n1109), .B2(new_n1104), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1097), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1100), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n965), .A2(new_n976), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1117), .A2(KEYINPUT121), .B1(new_n1026), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1120), .B(new_n1116), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n546), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(new_n546), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1110), .A2(new_n1115), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1108), .B1(new_n1126), .B2(KEYINPUT122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(KEYINPUT122), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1105), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1059), .A2(new_n962), .A3(new_n1061), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1073), .A2(new_n1133), .A3(new_n1065), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1074), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1070), .A2(G301), .A3(new_n1073), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1134), .B2(G171), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1058), .A2(new_n1136), .A3(new_n1084), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1093), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n966), .ZN(new_n1142));
  AND2_X1   g717(.A1(G290), .A2(G1986), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n984), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT110), .Z(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n979), .A3(new_n982), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n989), .B1(new_n1141), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g722(.A1(G227), .A2(new_n459), .ZN(new_n1149));
  AOI21_X1  g723(.A(new_n1149), .B1(new_n653), .B2(new_n655), .ZN(new_n1150));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1151));
  AND3_X1   g725(.A1(new_n1150), .A2(new_n1151), .A3(new_n697), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1150), .B2(new_n697), .ZN(new_n1153));
  OAI22_X1  g727(.A1(new_n897), .A2(new_n898), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g728(.A1(new_n959), .A2(new_n1154), .A3(KEYINPUT127), .ZN(new_n1155));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n1156));
  AND2_X1   g730(.A1(new_n895), .A2(new_n896), .ZN(new_n1157));
  INV_X1    g731(.A(new_n898), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n697), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n1159), .A2(KEYINPUT126), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n1150), .A2(new_n1151), .A3(new_n697), .ZN(new_n1161));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n947), .A2(new_n896), .ZN(new_n1163));
  OAI21_X1  g737(.A(KEYINPUT43), .B1(new_n1163), .B2(new_n951), .ZN(new_n1164));
  OR3_X1    g738(.A1(new_n951), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1156), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1155), .A2(new_n1167), .ZN(G308));
  OAI21_X1  g742(.A(KEYINPUT127), .B1(new_n959), .B2(new_n1154), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n1162), .A2(new_n1156), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1170), .ZN(G225));
endmodule


