//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n194), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n198), .A2(new_n200), .B1(KEYINPUT11), .B2(new_n195), .ZN(new_n207));
  NOR4_X1   g021(.A1(new_n207), .A2(G131), .A3(new_n204), .A4(new_n196), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(G128), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(G143), .B2(new_n211), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n217), .A3(G128), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT10), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT77), .A2(G104), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT78), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n227), .B(new_n228), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT79), .B(G101), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G107), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n231), .A2(KEYINPUT78), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n229), .A2(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n237), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n215), .B1(new_n218), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n221), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n248), .A3(new_n244), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n224), .A2(new_n245), .B1(new_n249), .B2(new_n223), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n254), .A3(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n215), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n220), .A2(KEYINPUT64), .A3(new_n257), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n212), .B2(new_n214), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n253), .A2(new_n255), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n250), .A2(new_n264), .A3(KEYINPUT81), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT81), .B1(new_n250), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n210), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n250), .A2(new_n264), .A3(new_n209), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n219), .A2(new_n221), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT80), .B(new_n249), .C1(new_n245), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n239), .B2(new_n244), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n201), .A2(new_n202), .ZN(new_n279));
  INV_X1    g093(.A(new_n196), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n205), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n279), .A2(new_n194), .A3(new_n280), .A4(new_n205), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n277), .A2(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n276), .A2(new_n284), .A3(KEYINPUT12), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT12), .B1(new_n276), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n268), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n272), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n267), .A2(new_n274), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n193), .B1(new_n289), .B2(G469), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n272), .B1(new_n267), .B2(new_n268), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n273), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n191), .B(new_n192), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n190), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G122), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT67), .A3(G116), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT2), .B(G113), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n253), .A2(new_n255), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n304), .A3(G116), .ZN(new_n312));
  OAI211_X1 g126(.A(G113), .B(new_n312), .C1(new_n306), .C2(new_n311), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n306), .A2(new_n307), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n245), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n309), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n310), .B1(new_n309), .B2(new_n316), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT6), .B(new_n299), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n255), .A2(new_n308), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT82), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n309), .A2(new_n310), .A3(new_n316), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n298), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n309), .A2(new_n298), .A3(new_n316), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT6), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n319), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n275), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n262), .A2(new_n261), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT64), .B1(new_n220), .B2(new_n257), .ZN(new_n333));
  AND4_X1   g147(.A1(KEYINPUT64), .A2(new_n212), .A3(new_n214), .A4(new_n257), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT83), .B(G224), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G953), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n329), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT7), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n343), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n298), .B(KEYINPUT8), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n245), .A2(new_n315), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n245), .A2(new_n315), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(KEYINPUT84), .B(new_n347), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n346), .A2(new_n352), .A3(new_n326), .A4(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n297), .B1(new_n341), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n299), .B1(new_n317), .B2(new_n318), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n327), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n357), .B2(new_n319), .ZN(new_n358));
  INV_X1    g172(.A(new_n297), .ZN(new_n359));
  INV_X1    g173(.A(new_n354), .ZN(new_n360));
  NOR4_X1   g174(.A1(new_n358), .A2(G902), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n295), .B(new_n296), .C1(new_n355), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n335), .B1(new_n282), .B2(new_n283), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n201), .A2(new_n195), .ZN(new_n365));
  NAND2_X1  g179(.A1(G134), .A2(G137), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(G131), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n283), .A2(new_n275), .A3(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n364), .A2(new_n368), .A3(new_n308), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n364), .C2(new_n368), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n263), .B1(new_n206), .B2(new_n208), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n283), .A2(new_n275), .A3(new_n367), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n369), .B1(new_n378), .B2(new_n308), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(G101), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G210), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n381), .B(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n308), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n371), .B2(new_n372), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT28), .B1(new_n369), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n371), .A2(new_n386), .A3(new_n372), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n192), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(G472), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n398));
  INV_X1    g212(.A(new_n384), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n308), .B1(new_n364), .B2(new_n368), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n400), .B2(new_n389), .ZN(new_n401));
  INV_X1    g215(.A(new_n391), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT31), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n403), .A2(new_n404), .B1(new_n379), .B2(new_n384), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n386), .B1(new_n370), .B2(new_n377), .ZN(new_n406));
  NOR4_X1   g220(.A1(new_n406), .A2(KEYINPUT31), .A3(new_n369), .A4(new_n399), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT69), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n373), .B(new_n374), .C1(new_n371), .C2(new_n372), .ZN(new_n409));
  AND4_X1   g223(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n376), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n308), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n389), .A3(new_n384), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n384), .B1(new_n388), .B2(new_n391), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(KEYINPUT31), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n379), .A2(new_n404), .A3(new_n384), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G472), .A2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n398), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT32), .B(new_n421), .C1(new_n408), .C2(new_n417), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n397), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G125), .B(G140), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT74), .B1(new_n424), .B2(new_n211), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n330), .A2(G140), .ZN(new_n426));
  INV_X1    g240(.A(G140), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G125), .ZN(new_n428));
  AND4_X1   g242(.A1(KEYINPUT74), .A2(new_n426), .A3(new_n428), .A4(new_n211), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n428), .A3(KEYINPUT72), .ZN(new_n430));
  OR3_X1    g244(.A1(new_n427), .A2(KEYINPUT72), .A3(G125), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n425), .A2(new_n429), .B1(new_n432), .B2(new_n211), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT18), .A2(G131), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n435));
  AOI21_X1  g249(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  INV_X1    g252(.A(G953), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(G214), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n213), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n441), .A2(KEYINPUT18), .A3(G131), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n430), .B2(new_n431), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n428), .A2(KEYINPUT16), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n211), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n448), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n427), .A2(KEYINPUT72), .A3(G125), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n424), .B2(KEYINPUT72), .ZN(new_n452));
  OAI211_X1 g266(.A(G146), .B(new_n450), .C1(new_n452), .C2(new_n446), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G131), .B1(new_n435), .B2(new_n436), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(new_n194), .A3(new_n442), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT17), .B(G131), .C1(new_n435), .C2(new_n436), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n445), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT86), .ZN(new_n463));
  OR2_X1    g277(.A1(G113), .A2(G122), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n465));
  NAND2_X1  g279(.A1(G113), .A2(G122), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n463), .A2(G104), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(G104), .B1(new_n463), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n461), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n445), .C1(new_n454), .C2(new_n460), .ZN(new_n473));
  AOI21_X1  g287(.A(G902), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT88), .B(G475), .Z(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT19), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT19), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n424), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n211), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n455), .A2(new_n457), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n453), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n477), .B(new_n470), .C1(new_n483), .C2(new_n445), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n445), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n471), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT20), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n473), .A2(KEYINPUT87), .B1(new_n471), .B2(new_n486), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(new_n489), .C1(new_n493), .C2(new_n484), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n476), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n439), .A2(G952), .ZN(new_n496));
  NAND2_X1  g310(.A1(G234), .A2(G237), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT92), .Z(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT21), .B(G898), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(G902), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT70), .B(G217), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n188), .A2(G953), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n213), .A2(G128), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n216), .B2(G143), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n201), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n230), .A2(new_n232), .ZN(new_n515));
  XOR2_X1   g329(.A(G116), .B(G122), .Z(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n216), .A2(G143), .ZN(new_n518));
  AND2_X1   g332(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n519));
  NOR2_X1   g333(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n520));
  OR3_X1    g334(.A1(new_n511), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n511), .B(new_n524), .C1(new_n519), .C2(new_n520), .ZN(new_n525));
  AND4_X1   g339(.A1(new_n518), .A2(new_n521), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n514), .B(new_n517), .C1(new_n526), .C2(new_n197), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n515), .A2(new_n516), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n301), .A2(KEYINPUT14), .A3(G122), .ZN(new_n529));
  OAI211_X1 g343(.A(G107), .B(new_n529), .C1(new_n516), .C2(KEYINPUT14), .ZN(new_n530));
  INV_X1    g344(.A(new_n514), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n513), .A2(new_n201), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n528), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n527), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n510), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n510), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n192), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G478), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n537), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n536), .B1(new_n527), .B2(new_n533), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n509), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  INV_X1    g362(.A(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n192), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n495), .A2(new_n506), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT93), .ZN(new_n552));
  AND2_X1   g366(.A1(KEYINPUT66), .A2(G128), .ZN(new_n553));
  NOR2_X1   g367(.A1(KEYINPUT66), .A2(G128), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT23), .B(G119), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n216), .A2(KEYINPUT71), .A3(KEYINPUT23), .A4(G119), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n304), .A2(G128), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT23), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n304), .B2(G128), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n216), .A2(G119), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(new_n559), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  OAI22_X1  g379(.A1(new_n562), .A2(G110), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n453), .C1(new_n425), .C2(new_n429), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n563), .A2(new_n559), .A3(new_n565), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n449), .B2(new_n453), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(G110), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(KEYINPUT73), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT73), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT75), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n439), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT22), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n195), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n567), .C1(new_n571), .C2(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n192), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n508), .B1(G234), .B2(new_n192), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n588), .A3(new_n192), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n587), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n363), .A2(new_n423), .A3(new_n552), .A4(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(new_n234), .Z(G3));
  NOR3_X1   g410(.A1(new_n405), .A2(KEYINPUT69), .A3(new_n407), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n419), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n408), .B2(new_n417), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n295), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n593), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n506), .B(new_n296), .C1(new_n361), .C2(new_n355), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n534), .A2(KEYINPUT94), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n509), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n510), .B1(new_n534), .B2(KEYINPUT94), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(KEYINPUT33), .B2(new_n548), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(G478), .A3(new_n192), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n541), .A2(new_n542), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n495), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  AOI21_X1  g431(.A(new_n549), .B1(new_n548), .B2(new_n192), .ZN(new_n618));
  AOI211_X1 g432(.A(G902), .B(new_n543), .C1(new_n547), .C2(new_n539), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n476), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n491), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n491), .B2(new_n494), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n604), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n603), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  INV_X1    g445(.A(KEYINPUT93), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n551), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n362), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n588), .B1(new_n584), .B2(new_n192), .ZN(new_n635));
  AOI211_X1 g449(.A(KEYINPUT25), .B(G902), .C1(new_n582), .C2(new_n583), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n574), .A2(new_n581), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n579), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n637), .A2(new_n587), .B1(new_n591), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G110), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  NAND2_X1  g461(.A1(new_n599), .A2(KEYINPUT32), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n421), .B1(new_n408), .B2(new_n417), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n398), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n641), .B1(new_n651), .B2(new_n397), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n500), .B1(new_n653), .B2(new_n504), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n626), .A2(new_n621), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n329), .A2(new_n340), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n354), .A3(new_n192), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n359), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n341), .A2(new_n297), .A3(new_n354), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n657), .A2(new_n662), .A3(KEYINPUT97), .A4(new_n296), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n296), .B1(new_n361), .B2(new_n355), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n656), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n652), .A2(new_n663), .A3(new_n295), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n246), .ZN(G30));
  NAND2_X1  g483(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n660), .A2(new_n671), .A3(new_n661), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT38), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(KEYINPUT38), .A3(new_n672), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n379), .A2(new_n399), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n400), .A2(new_n389), .A3(new_n399), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n192), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n651), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n640), .A2(new_n591), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n590), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n495), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n544), .A2(new_n550), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n676), .A2(KEYINPUT100), .A3(new_n296), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n675), .A3(new_n674), .A4(new_n296), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n654), .B(KEYINPUT101), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n295), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  NAND3_X1  g510(.A1(new_n689), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n692), .A3(new_n699), .A4(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n213), .ZN(G45));
  NOR2_X1   g516(.A1(new_n613), .A2(new_n654), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n652), .A2(new_n363), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  OAI21_X1  g519(.A(new_n192), .B1(new_n291), .B2(new_n293), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n189), .A3(new_n294), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n614), .A2(new_n423), .A3(new_n594), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n628), .A2(new_n423), .A3(new_n594), .A4(new_n709), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n665), .A2(new_n708), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n423), .A3(new_n552), .A4(new_n683), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n421), .B1(new_n405), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n414), .A2(KEYINPUT104), .A3(new_n416), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n724));
  OAI22_X1  g538(.A1(new_n723), .A2(new_n724), .B1(new_n600), .B2(new_n601), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n593), .ZN(new_n726));
  INV_X1    g540(.A(new_n686), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n506), .A3(new_n715), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT106), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(G122), .Z(G24));
  NOR2_X1   g544(.A1(new_n725), .A2(new_n641), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n703), .A3(new_n715), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND3_X1  g547(.A1(new_n660), .A2(new_n296), .A3(new_n661), .ZN(new_n734));
  INV_X1    g548(.A(new_n295), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n423), .A2(new_n736), .A3(new_n594), .A4(new_n703), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n593), .B1(new_n651), .B2(new_n397), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n703), .A4(new_n736), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  AND3_X1   g557(.A1(new_n740), .A2(new_n657), .A3(new_n736), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n197), .ZN(G36));
  OR2_X1    g559(.A1(new_n289), .A2(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n289), .A2(KEYINPUT45), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(G469), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n193), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n748), .B2(new_n749), .ZN(new_n753));
  INV_X1    g567(.A(new_n294), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n190), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n694), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n610), .A2(new_n611), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n495), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT43), .A3(new_n495), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n642), .A3(new_n683), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n734), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n758), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT108), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(new_n703), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n753), .A2(new_n754), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n189), .B1(new_n775), .B2(new_n752), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n773), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n734), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n423), .A2(new_n594), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n779), .A2(KEYINPUT109), .A3(new_n780), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n707), .A2(new_n294), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n594), .B(new_n296), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n190), .A3(new_n760), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT110), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n674), .A2(new_n675), .ZN(new_n794));
  INV_X1    g608(.A(new_n681), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n790), .A2(new_n788), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n774), .B(new_n778), .C1(new_n189), .C2(new_n789), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n499), .B1(new_n762), .B2(new_n763), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n726), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n780), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT51), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n734), .A2(new_n708), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n799), .A2(new_n731), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n708), .A2(new_n296), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT116), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n794), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n810), .B2(new_n811), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n802), .B(new_n807), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n795), .A2(new_n500), .A3(new_n594), .A4(new_n806), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n759), .A2(new_n684), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n805), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n802), .A2(new_n807), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n802), .B2(new_n803), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n814), .A2(new_n815), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n825), .A3(new_n826), .A4(new_n820), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n822), .A2(new_n827), .A3(new_n496), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n818), .A2(new_n612), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n710), .A2(new_n728), .A3(new_n713), .A4(new_n716), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n634), .B1(new_n740), .B2(new_n643), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n620), .A2(new_n684), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n612), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n604), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n603), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT111), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(KEYINPUT111), .A2(new_n595), .A3(new_n644), .A4(new_n836), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n744), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n731), .A2(new_n703), .A3(new_n736), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n734), .A2(new_n735), .A3(new_n476), .A4(new_n654), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n652), .A2(new_n842), .A3(new_n620), .A4(new_n626), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n742), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n830), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n728), .A2(new_n710), .A3(new_n713), .A4(new_n716), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n552), .A2(new_n296), .A3(new_n662), .A4(new_n295), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n423), .A2(new_n594), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n683), .B(new_n599), .C1(new_n601), .C2(new_n600), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n836), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n832), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n744), .B1(new_n739), .B2(new_n741), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n843), .A2(new_n841), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(KEYINPUT112), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n845), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n654), .B(KEYINPUT113), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n681), .A2(new_n363), .A3(new_n687), .A4(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n667), .A2(new_n704), .A3(new_n732), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n864));
  OAI21_X1  g678(.A(KEYINPUT115), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n667), .A2(new_n704), .A3(new_n732), .A4(new_n862), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  INV_X1    g682(.A(new_n864), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n859), .A2(new_n860), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n845), .A2(new_n858), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n872), .B(KEYINPUT54), .C1(new_n860), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n839), .A2(new_n844), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n876), .B(new_n878), .C1(new_n874), .C2(KEYINPUT53), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n828), .A2(new_n829), .A3(new_n875), .A4(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n800), .A2(new_n665), .A3(new_n708), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n740), .A2(new_n799), .A3(new_n806), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  NOR3_X1   g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n797), .B1(new_n884), .B2(new_n885), .ZN(G75));
  XNOR2_X1  g700(.A(new_n329), .B(new_n339), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n873), .A2(new_n866), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n859), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n871), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n891));
  OAI211_X1 g705(.A(G210), .B(G902), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT55), .ZN(new_n893));
  NOR2_X1   g707(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT55), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n887), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n439), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n897), .A2(new_n901), .A3(new_n903), .ZN(G51));
  OAI21_X1  g718(.A(new_n878), .B1(new_n874), .B2(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n879), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n909), .A2(new_n910), .B1(new_n291), .B2(new_n293), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n905), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n748), .B(KEYINPUT120), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n902), .B1(new_n911), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n912), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n488), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n488), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n902), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n906), .B2(new_n879), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n609), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT122), .B1(new_n925), .B2(new_n609), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n875), .B2(new_n879), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n903), .B1(new_n928), .B2(new_n609), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n905), .A2(new_n640), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n905), .A2(KEYINPUT123), .A3(new_n640), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n905), .A2(new_n933), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n584), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n584), .B1(new_n905), .B2(new_n933), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(KEYINPUT124), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n938), .A2(new_n941), .A3(new_n944), .A4(new_n903), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n902), .B(new_n943), .C1(new_n936), .C2(new_n937), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(KEYINPUT61), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n502), .B2(new_n337), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n855), .B2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n357), .B(new_n319), .C1(G898), .C2(new_n439), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  OAI21_X1  g766(.A(G953), .B1(new_n270), .B2(new_n653), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n439), .A2(G900), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n478), .A2(new_n480), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n378), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n786), .A2(new_n770), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n667), .A2(new_n704), .A3(new_n732), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n665), .A2(new_n686), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n758), .A2(new_n740), .A3(new_n769), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n958), .A2(new_n960), .A3(new_n856), .A4(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n954), .B(new_n957), .C1(new_n963), .C2(new_n439), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n701), .B2(new_n959), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n698), .A2(KEYINPUT62), .A3(new_n700), .A4(new_n960), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n612), .A2(new_n833), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n740), .A2(new_n694), .A3(new_n736), .A4(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n971), .A2(new_n439), .A3(new_n957), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n953), .B1(new_n964), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n963), .A2(new_n439), .ZN(new_n974));
  INV_X1    g788(.A(new_n954), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n956), .ZN(new_n976));
  INV_X1    g790(.A(new_n953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n971), .A2(new_n439), .A3(new_n957), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n973), .A2(new_n979), .ZN(G72));
  NAND4_X1  g794(.A1(new_n968), .A2(new_n958), .A3(new_n855), .A4(new_n970), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n601), .A2(new_n192), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n902), .B1(new_n985), .B2(new_n677), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n859), .A2(new_n889), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n871), .A2(new_n860), .ZN(new_n988));
  AOI22_X1  g802(.A1(KEYINPUT53), .A2(new_n987), .B1(new_n988), .B2(new_n859), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n406), .A2(new_n369), .A3(new_n384), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n677), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n984), .A4(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n984), .B1(new_n963), .B2(new_n839), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n990), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n986), .A2(new_n996), .A3(new_n998), .ZN(G57));
endmodule


