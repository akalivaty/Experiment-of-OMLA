

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XNOR2_X1 U326 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U327 ( .A(n439), .B(n438), .ZN(n471) );
  XOR2_X1 U328 ( .A(KEYINPUT41), .B(n581), .Z(n571) );
  XOR2_X1 U329 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n294) );
  XOR2_X1 U330 ( .A(KEYINPUT13), .B(G57GAT), .Z(n295) );
  XOR2_X1 U331 ( .A(n381), .B(n336), .Z(n296) );
  AND2_X1 U332 ( .A1(n474), .A2(n473), .ZN(n297) );
  INV_X1 U333 ( .A(KEYINPUT10), .ZN(n338) );
  INV_X1 U334 ( .A(n523), .ZN(n473) );
  NOR2_X1 U335 ( .A1(n451), .A2(n450), .ZN(n490) );
  XNOR2_X1 U336 ( .A(n341), .B(n340), .ZN(n345) );
  NOR2_X1 U337 ( .A1(n591), .A2(n453), .ZN(n454) );
  XOR2_X1 U338 ( .A(KEYINPUT48), .B(n470), .Z(n553) );
  OR2_X1 U339 ( .A1(n492), .A2(n522), .ZN(n455) );
  XOR2_X1 U340 ( .A(n429), .B(n426), .Z(n537) );
  XNOR2_X1 U341 ( .A(n481), .B(G190GAT), .ZN(n482) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n456) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n299) );
  NAND2_X1 U346 ( .A1(G230GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n300), .B(KEYINPUT71), .Z(n305) );
  XOR2_X1 U349 ( .A(G92GAT), .B(G85GAT), .Z(n302) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n347) );
  XNOR2_X1 U352 ( .A(G71GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n295), .B(n303), .ZN(n360) );
  XNOR2_X1 U354 ( .A(n347), .B(n360), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U356 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n307) );
  XNOR2_X1 U357 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U359 ( .A(n309), .B(n308), .Z(n311) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G148GAT), .Z(n397) );
  XOR2_X1 U361 ( .A(G176GAT), .B(G64GAT), .Z(n430) );
  XNOR2_X1 U362 ( .A(n397), .B(n430), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n581) );
  XOR2_X1 U364 ( .A(KEYINPUT66), .B(G8GAT), .Z(n313) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n334) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n315) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G197GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U370 ( .A(G36GAT), .B(G50GAT), .Z(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n330) );
  XNOR2_X1 U372 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n318), .B(KEYINPUT70), .ZN(n319) );
  XOR2_X1 U374 ( .A(n319), .B(KEYINPUT29), .Z(n328) );
  INV_X1 U375 ( .A(G43GAT), .ZN(n320) );
  NAND2_X1 U376 ( .A1(G29GAT), .A2(n320), .ZN(n323) );
  INV_X1 U377 ( .A(G29GAT), .ZN(n321) );
  NAND2_X1 U378 ( .A1(n321), .A2(G43GAT), .ZN(n322) );
  NAND2_X1 U379 ( .A1(n323), .A2(n322), .ZN(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n336) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n326), .B(KEYINPUT68), .ZN(n357) );
  XNOR2_X1 U384 ( .A(n336), .B(n357), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n332) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n565) );
  INV_X1 U390 ( .A(n565), .ZN(n576) );
  NOR2_X1 U391 ( .A1(n581), .A2(n576), .ZN(n335) );
  XOR2_X1 U392 ( .A(n335), .B(KEYINPUT74), .Z(n492) );
  XNOR2_X1 U393 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n350) );
  XOR2_X1 U394 ( .A(G134GAT), .B(KEYINPUT76), .Z(n381) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n296), .B(n337), .ZN(n341) );
  XOR2_X1 U397 ( .A(G50GAT), .B(G162GAT), .Z(n401) );
  XNOR2_X1 U398 ( .A(n401), .B(KEYINPUT77), .ZN(n339) );
  XOR2_X1 U399 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n343) );
  XNOR2_X1 U400 ( .A(KEYINPUT9), .B(KEYINPUT75), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U402 ( .A(n345), .B(n344), .Z(n349) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n346), .B(G218GAT), .ZN(n435) );
  XNOR2_X1 U405 ( .A(n435), .B(n347), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n562) );
  XNOR2_X1 U407 ( .A(n562), .B(KEYINPUT78), .ZN(n480) );
  XNOR2_X1 U408 ( .A(n350), .B(n480), .ZN(n591) );
  XOR2_X1 U409 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n352) );
  XNOR2_X1 U410 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U412 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n354) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U415 ( .A(n355), .B(KEYINPUT79), .Z(n359) );
  XOR2_X1 U416 ( .A(G8GAT), .B(G183GAT), .Z(n356) );
  XOR2_X1 U417 ( .A(G211GAT), .B(n356), .Z(n427) );
  XNOR2_X1 U418 ( .A(n357), .B(n427), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n361) );
  XOR2_X1 U420 ( .A(n361), .B(n360), .Z(n363) );
  XOR2_X1 U421 ( .A(G15GAT), .B(G127GAT), .Z(n414) );
  XOR2_X1 U422 ( .A(G22GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U423 ( .A(n414), .B(n396), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U425 ( .A(n365), .B(n364), .Z(n560) );
  XOR2_X1 U426 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n367) );
  XNOR2_X1 U427 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U429 ( .A(G141GAT), .B(n368), .Z(n409) );
  XOR2_X1 U430 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n370) );
  XNOR2_X1 U431 ( .A(G1GAT), .B(G57GAT), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U433 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n372) );
  XNOR2_X1 U434 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U436 ( .A(n374), .B(n373), .Z(n388) );
  XOR2_X1 U437 ( .A(G120GAT), .B(KEYINPUT82), .Z(n376) );
  XNOR2_X1 U438 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n413) );
  XOR2_X1 U440 ( .A(n413), .B(KEYINPUT92), .Z(n378) );
  NAND2_X1 U441 ( .A1(G225GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U443 ( .A(G85GAT), .B(G155GAT), .Z(n380) );
  XNOR2_X1 U444 ( .A(G127GAT), .B(G162GAT), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U446 ( .A(n382), .B(n381), .Z(n384) );
  XNOR2_X1 U447 ( .A(G29GAT), .B(G148GAT), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n409), .B(n389), .ZN(n523) );
  XOR2_X1 U452 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n391) );
  XNOR2_X1 U453 ( .A(G218GAT), .B(G106GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U455 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n393) );
  XNOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT24), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n395), .B(n394), .Z(n403) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U460 ( .A1(G228GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U464 ( .A(n404), .B(G78GAT), .Z(n407) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n405), .B(KEYINPUT21), .ZN(n428) );
  XNOR2_X1 U467 ( .A(n428), .B(KEYINPUT86), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n475) );
  INV_X1 U470 ( .A(n475), .ZN(n441) );
  XNOR2_X1 U471 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n294), .B(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n429) );
  XOR2_X1 U475 ( .A(n414), .B(n413), .Z(n416) );
  XNOR2_X1 U476 ( .A(G190GAT), .B(G99GAT), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U478 ( .A(G183GAT), .B(G176GAT), .Z(n418) );
  NAND2_X1 U479 ( .A1(G227GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n420), .B(n419), .Z(n425) );
  XOR2_X1 U482 ( .A(KEYINPUT83), .B(G71GAT), .Z(n422) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G134GAT), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n423), .B(KEYINPUT20), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U487 ( .A(n537), .ZN(n479) );
  XOR2_X1 U488 ( .A(n428), .B(n427), .Z(n439) );
  INV_X1 U489 ( .A(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U493 ( .A(n434), .B(G92GAT), .Z(n437) );
  XNOR2_X1 U494 ( .A(G204GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  NOR2_X1 U496 ( .A1(n479), .A2(n471), .ZN(n440) );
  NOR2_X1 U497 ( .A1(n441), .A2(n440), .ZN(n442) );
  XOR2_X1 U498 ( .A(KEYINPUT25), .B(n442), .Z(n445) );
  NOR2_X1 U499 ( .A1(n537), .A2(n475), .ZN(n443) );
  XNOR2_X1 U500 ( .A(KEYINPUT26), .B(n443), .ZN(n575) );
  INV_X1 U501 ( .A(n471), .ZN(n526) );
  XNOR2_X1 U502 ( .A(KEYINPUT27), .B(n526), .ZN(n447) );
  AND2_X1 U503 ( .A1(n575), .A2(n447), .ZN(n444) );
  NOR2_X1 U504 ( .A1(n445), .A2(n444), .ZN(n446) );
  NOR2_X1 U505 ( .A1(n523), .A2(n446), .ZN(n451) );
  NAND2_X1 U506 ( .A1(n447), .A2(n523), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n448), .B(KEYINPUT95), .ZN(n551) );
  XOR2_X1 U508 ( .A(KEYINPUT28), .B(n475), .Z(n530) );
  INV_X1 U509 ( .A(n530), .ZN(n449) );
  NAND2_X1 U510 ( .A1(n551), .A2(n449), .ZN(n536) );
  NOR2_X1 U511 ( .A1(n536), .A2(n537), .ZN(n450) );
  NOR2_X1 U512 ( .A1(n560), .A2(n490), .ZN(n452) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(n452), .Z(n453) );
  XNOR2_X1 U514 ( .A(KEYINPUT37), .B(n454), .ZN(n522) );
  XOR2_X1 U515 ( .A(KEYINPUT38), .B(n455), .Z(n509) );
  NAND2_X1 U516 ( .A1(n509), .A2(n537), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT111), .B(n560), .ZN(n544) );
  XOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n459) );
  NAND2_X1 U519 ( .A1(n571), .A2(n565), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n562), .A2(n460), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n544), .A2(n461), .ZN(n462) );
  XNOR2_X1 U523 ( .A(KEYINPUT47), .B(n462), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT113), .ZN(n469) );
  INV_X1 U525 ( .A(n560), .ZN(n587) );
  NOR2_X1 U526 ( .A1(n587), .A2(n591), .ZN(n465) );
  XNOR2_X1 U527 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U529 ( .A1(n466), .A2(n581), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n576), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n471), .A2(n553), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT54), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n297), .A2(n475), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X2 U537 ( .A1(n479), .A2(n478), .ZN(n572) );
  NAND2_X1 U538 ( .A1(n572), .A2(n480), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n481) );
  INV_X1 U540 ( .A(n572), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n484), .A2(n544), .ZN(n487) );
  INV_X1 U542 ( .A(G183GAT), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n485), .B(KEYINPUT122), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1350GAT) );
  NOR2_X1 U545 ( .A1(n587), .A2(n480), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  NOR2_X1 U547 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U548 ( .A(KEYINPUT96), .B(n491), .Z(n511) );
  NOR2_X1 U549 ( .A1(n492), .A2(n511), .ZN(n501) );
  NAND2_X1 U550 ( .A1(n523), .A2(n501), .ZN(n496) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n494) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n501), .A2(n526), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n499) );
  NAND2_X1 U558 ( .A1(n501), .A2(n537), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U560 ( .A(G15GAT), .B(n500), .Z(G1326GAT) );
  NAND2_X1 U561 ( .A1(n530), .A2(n501), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  NAND2_X1 U564 ( .A1(n509), .A2(n523), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT103), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n526), .A2(n509), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n530), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n514) );
  NAND2_X1 U574 ( .A1(n576), .A2(n571), .ZN(n521) );
  NOR2_X1 U575 ( .A1(n521), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT106), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n518), .A2(n523), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n526), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n537), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n530), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT107), .Z(n525) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n531), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT108), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n537), .A2(n531), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n535) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n533) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n553), .A2(n536), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n576), .A2(n543), .ZN(n539) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  INV_X1 U605 ( .A(n543), .ZN(n547) );
  AND2_X1 U606 ( .A1(n571), .A2(n547), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n480), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n575), .ZN(n552) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n565), .A2(n563), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(n557), .Z(n559) );
  NAND2_X1 U625 ( .A1(n563), .A2(n571), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT119), .Z(n567) );
  NAND2_X1 U632 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT120), .B(n570), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n297), .A2(n575), .ZN(n590) );
  NOR2_X1 U641 ( .A1(n576), .A2(n590), .ZN(n580) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT124), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n590), .A2(n582), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U652 ( .A1(n587), .A2(n590), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

