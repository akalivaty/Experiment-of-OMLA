//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n188), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT67), .A3(G137), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n189), .A2(new_n191), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n190), .B2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n190), .A2(G137), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n196), .A2(KEYINPUT71), .A3(new_n202), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G143), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n211), .A2(new_n212), .B1(KEYINPUT1), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n205), .A2(new_n206), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n210), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n221), .B(new_n222), .C1(new_n225), .C2(new_n215), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n209), .A2(G146), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n228), .A2(new_n213), .B1(new_n224), .B2(new_n223), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n222), .B1(new_n229), .B2(new_n221), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n198), .A2(new_n201), .A3(new_n199), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n202), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(KEYINPUT30), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(G119), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT69), .A4(G119), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(G119), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT2), .B(G113), .Z(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n243), .A2(new_n248), .A3(new_n244), .A4(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n229), .A2(new_n221), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n229), .A2(new_n255), .A3(new_n221), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n234), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n218), .A2(new_n202), .A3(new_n196), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n236), .A2(new_n252), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n252), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n219), .A2(new_n263), .A3(new_n235), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n267), .B(KEYINPUT27), .Z(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT26), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(G101), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT31), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n264), .A2(new_n272), .B1(new_n252), .B2(new_n259), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n219), .A2(new_n263), .A3(KEYINPUT28), .A4(new_n235), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  INV_X1    g090(.A(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n269), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n262), .A3(new_n279), .A4(new_n264), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(KEYINPUT32), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n265), .A2(new_n278), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n263), .B1(new_n219), .B2(new_n235), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n264), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT72), .B(new_n263), .C1(new_n235), .C2(new_n219), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT28), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n264), .A2(new_n272), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(KEYINPUT29), .A3(new_n278), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n288), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n281), .A2(new_n299), .A3(KEYINPUT32), .A4(new_n282), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n281), .A2(new_n282), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n284), .A2(new_n298), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT77), .B(G125), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT16), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G125), .A2(G140), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n305), .B2(G140), .ZN(new_n310));
  OAI211_X1 g124(.A(G146), .B(new_n308), .C1(new_n310), .C2(new_n306), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n207), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n212), .A2(G119), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT78), .B1(new_n322), .B2(G110), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n319), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(KEYINPUT75), .B2(new_n318), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n322), .A2(KEYINPUT78), .A3(G110), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n311), .B(new_n313), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n326), .A2(new_n328), .B1(G110), .B2(new_n322), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT77), .A2(G125), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT77), .A2(G125), .ZN(new_n334));
  OAI21_X1  g148(.A(G140), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n309), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n306), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n306), .A2(new_n307), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n207), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n311), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(G221), .A3(G234), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT22), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n331), .A2(new_n343), .A3(new_n348), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G217), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(G234), .B2(new_n296), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(G902), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n356), .A2(KEYINPUT79), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n296), .A3(new_n351), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT25), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n354), .B(KEYINPUT74), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n358), .B2(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(KEYINPUT79), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n304), .A2(KEYINPUT80), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT80), .B1(new_n304), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G214), .B1(G237), .B2(G902), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G101), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(KEYINPUT82), .A3(new_n377), .A4(G101), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n371), .A2(new_n374), .A3(new_n277), .A4(new_n375), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n377), .B1(new_n376), .B2(G101), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n252), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n244), .A4(new_n246), .ZN(new_n386));
  INV_X1    g200(.A(G113), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n245), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n370), .A2(G107), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n373), .A2(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n382), .A2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT83), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n390), .A2(new_n396), .A3(new_n251), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT86), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT88), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n407), .A3(new_n401), .A4(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n401), .B1(new_n400), .B2(new_n404), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n396), .A2(new_n398), .ZN(new_n412));
  INV_X1    g226(.A(new_n247), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n413), .A2(new_n248), .B1(new_n386), .B2(new_n389), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n412), .A2(new_n414), .B1(new_n384), .B2(new_n252), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n415), .B2(new_n403), .ZN(new_n416));
  AND4_X1   g230(.A1(new_n411), .A2(new_n385), .A3(new_n399), .A4(new_n403), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n410), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n214), .A2(new_n217), .A3(new_n338), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n229), .A2(new_n221), .A3(new_n305), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G224), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n421), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n409), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n420), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  OAI22_X1  g243(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(new_n423), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n431), .A2(KEYINPUT90), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n431), .B2(KEYINPUT90), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n419), .A2(new_n420), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n414), .A2(new_n397), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n414), .A2(new_n397), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n403), .B(KEYINPUT8), .Z(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT87), .B1(new_n400), .B2(new_n404), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n415), .A2(new_n411), .A3(new_n403), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n425), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n425), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n369), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT92), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n209), .A2(G128), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT96), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n212), .A2(G143), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n452), .A2(KEYINPUT96), .A3(new_n453), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT13), .B1(new_n209), .B2(G128), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT95), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n190), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT97), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT97), .B1(new_n452), .B2(new_n455), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n190), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n238), .A2(new_n240), .A3(G122), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n237), .A2(G122), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n465), .A2(new_n373), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n373), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n455), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT97), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(G134), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n467), .B1(new_n464), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n465), .A2(new_n478), .A3(new_n466), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT14), .A4(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G107), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n479), .A2(KEYINPUT98), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n480), .A2(G107), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n465), .A2(new_n478), .A3(new_n466), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT99), .B(new_n477), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT98), .B1(new_n479), .B2(new_n481), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n483), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT99), .B1(new_n491), .B2(new_n477), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n471), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT9), .B(G234), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(new_n353), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n477), .B1(new_n482), .B2(new_n486), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT99), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n487), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n471), .A3(new_n495), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  OAI22_X1  g318(.A1(new_n503), .A2(KEYINPUT100), .B1(KEYINPUT15), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n495), .B1(new_n501), .B2(new_n471), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n470), .B(new_n496), .C1(new_n500), .C2(new_n487), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n296), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT100), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n503), .A2(KEYINPUT100), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G113), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(new_n370), .ZN(new_n516));
  INV_X1    g330(.A(G237), .ZN(new_n517));
  AND4_X1   g331(.A1(G143), .A2(new_n517), .A3(new_n345), .A4(G214), .ZN(new_n518));
  AOI21_X1  g332(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n345), .A3(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n209), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n200), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT17), .B(G131), .C1(new_n518), .C2(new_n519), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n341), .A2(new_n311), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n335), .A2(new_n336), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n313), .B1(new_n529), .B2(new_n207), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n524), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT18), .B(G131), .C1(new_n518), .C2(new_n519), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n516), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n516), .B(new_n534), .C1(new_n342), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n528), .A2(KEYINPUT93), .A3(new_n516), .A4(new_n534), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G475), .B1(new_n541), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n520), .A2(new_n525), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n312), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n529), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n311), .B(new_n545), .C1(new_n548), .C2(G146), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n516), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n550), .B1(new_n539), .B2(new_n540), .ZN(new_n559));
  INV_X1    g373(.A(new_n554), .ZN(new_n560));
  NOR4_X1   g374(.A1(new_n559), .A2(new_n557), .A3(KEYINPUT20), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n543), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n514), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n565), .A2(G952), .A3(new_n345), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n345), .A2(G227), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n234), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n218), .A2(new_n394), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n397), .A2(new_n217), .A3(new_n214), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n380), .A2(new_n381), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n383), .A2(new_n382), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n231), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n396), .A2(KEYINPUT10), .A3(new_n218), .A4(new_n398), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n583), .A2(new_n575), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n574), .B1(new_n580), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n586), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n234), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n574), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n571), .B1(new_n595), .B2(new_n296), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n587), .A2(KEYINPUT84), .A3(new_n593), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT84), .B1(new_n587), .B2(new_n593), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n597), .A2(new_n598), .A3(new_n580), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n592), .B2(new_n587), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n571), .B(new_n296), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n593), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n578), .B(KEYINPUT12), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n587), .A2(KEYINPUT84), .A3(new_n593), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n600), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT85), .A3(new_n571), .A4(new_n296), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n596), .B1(new_n603), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G221), .B1(new_n494), .B2(G902), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT81), .Z(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n451), .A2(new_n570), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n368), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n277), .ZN(G3));
  AND3_X1   g433(.A1(new_n425), .A2(new_n444), .A3(new_n446), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n446), .B1(new_n425), .B2(new_n444), .ZN(new_n621));
  INV_X1    g435(.A(new_n369), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n569), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(KEYINPUT94), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n542), .B1(new_n628), .B2(new_n561), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n506), .B2(new_n507), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n497), .A2(KEYINPUT33), .A3(new_n502), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n504), .A2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n508), .A2(new_n504), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n281), .B2(new_n296), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n301), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n613), .A3(new_n615), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n638), .A2(new_n365), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  OAI21_X1  g460(.A(new_n542), .B1(new_n556), .B2(new_n626), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n625), .A2(new_n514), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n365), .A3(new_n643), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n344), .B(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n359), .A2(new_n361), .B1(new_n355), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n451), .A2(new_n643), .A3(new_n570), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AND3_X1   g472(.A1(new_n616), .A2(new_n304), .A3(new_n655), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  INV_X1    g474(.A(new_n566), .ZN(new_n661));
  INV_X1    g475(.A(new_n567), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(G900), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n542), .B(new_n663), .C1(new_n556), .C2(new_n626), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n623), .A2(new_n660), .A3(new_n513), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n425), .A2(new_n444), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n445), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n425), .A2(new_n444), .A3(new_n446), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n369), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n513), .A2(new_n665), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT101), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n659), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XNOR2_X1  g489(.A(new_n663), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n616), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n265), .A2(new_n278), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n291), .A2(new_n292), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n681), .B(new_n296), .C1(new_n682), .C2(new_n278), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G472), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n284), .A2(new_n303), .A3(new_n300), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(new_n448), .B2(new_n449), .ZN(new_n688));
  INV_X1    g502(.A(new_n447), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n667), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n425), .A2(new_n444), .A3(new_n447), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(KEYINPUT38), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n629), .A2(new_n513), .A3(new_n369), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n686), .A2(new_n693), .A3(new_n655), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n679), .A2(new_n680), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT103), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  NAND3_X1  g512(.A1(new_n629), .A2(new_n636), .A3(new_n663), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n670), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n616), .A3(new_n304), .A4(new_n655), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  AND2_X1   g516(.A1(new_n304), .A2(new_n365), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n603), .A2(new_n612), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n571), .B1(new_n611), .B2(new_n296), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n704), .A2(new_n614), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(new_n614), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n709), .B(new_n705), .C1(new_n603), .C2(new_n612), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n703), .A2(new_n638), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n648), .A2(new_n703), .A3(new_n708), .A4(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NOR2_X1   g531(.A1(new_n707), .A2(new_n670), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n304), .A3(new_n570), .A4(new_n655), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NOR4_X1   g534(.A1(new_n670), .A2(new_n514), .A3(new_n563), .A4(new_n569), .ZN(new_n721));
  INV_X1    g535(.A(new_n282), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n293), .A2(new_n294), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n270), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n271), .A2(new_n280), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n364), .A2(new_n640), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n712), .A3(new_n727), .A4(new_n708), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NOR3_X1   g543(.A1(new_n726), .A2(new_n654), .A3(new_n640), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n629), .A2(new_n732), .A3(new_n636), .A4(new_n663), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n718), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n613), .A2(new_n709), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n690), .A2(new_n369), .A3(new_n691), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n304), .A3(new_n365), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n731), .A2(new_n733), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n736), .C1(new_n740), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n303), .A2(KEYINPUT107), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n303), .A2(KEYINPUT107), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n283), .A3(new_n298), .A4(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n365), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n741), .A2(new_n736), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n737), .A3(new_n739), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  OR2_X1    g568(.A1(new_n740), .A2(new_n671), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  AND2_X1   g570(.A1(new_n634), .A2(new_n635), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n629), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n636), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n634), .A2(new_n762), .A3(new_n635), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n563), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n642), .A2(new_n758), .A3(new_n764), .A4(new_n655), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT44), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  INV_X1    g581(.A(new_n591), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n575), .B1(new_n768), .B2(new_n583), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n604), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n593), .B1(new_n607), .B2(new_n587), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n589), .A2(KEYINPUT45), .A3(new_n594), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(G469), .ZN(new_n774));
  NAND2_X1  g588(.A1(G469), .A2(G902), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT46), .B1(new_n774), .B2(new_n775), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n603), .B2(new_n612), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n781), .A2(new_n614), .A3(new_n676), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n738), .B(KEYINPUT110), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n766), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n781), .B2(new_n614), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n709), .B(new_n789), .C1(new_n778), .C2(new_n780), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n304), .A2(new_n365), .A3(new_n699), .A4(new_n738), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT112), .Z(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n307), .ZN(G42));
  NOR2_X1   g609(.A1(new_n707), .A2(new_n738), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n365), .A3(new_n566), .A4(new_n686), .ZN(new_n797));
  OAI211_X1 g611(.A(G952), .B(new_n345), .C1(new_n797), .C2(new_n637), .ZN(new_n798));
  INV_X1    g612(.A(new_n727), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n758), .A2(new_n764), .A3(new_n566), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n758), .A2(new_n764), .A3(new_n802), .A4(new_n566), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n798), .B1(new_n718), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n803), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n796), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT48), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n750), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n807), .B2(new_n750), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n797), .A2(new_n629), .A3(new_n636), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n807), .B2(new_n730), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n705), .B1(new_n603), .B2(new_n612), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n615), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n788), .B2(new_n790), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n783), .A3(new_n804), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n369), .B1(new_n688), .B2(new_n692), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n710), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n822), .A3(new_n710), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT50), .A3(new_n804), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n804), .A3(KEYINPUT118), .A4(KEYINPUT50), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n804), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n833), .B(KEYINPUT50), .C1(new_n824), .C2(new_n804), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n818), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n811), .B1(new_n836), .B2(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n806), .A2(new_n727), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n822), .A2(new_n710), .A3(new_n693), .A4(new_n622), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n822), .B1(new_n819), .B2(new_n710), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n831), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n833), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n830), .A2(KEYINPUT117), .A3(new_n831), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n827), .A3(new_n828), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n813), .A2(new_n817), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n850), .B(KEYINPUT51), .C1(new_n845), .C2(new_n846), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n837), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n668), .A2(new_n669), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n694), .A2(new_n613), .A3(new_n855), .A4(new_n709), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n654), .A2(new_n663), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n685), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n659), .A2(new_n673), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT113), .A3(new_n701), .A4(new_n734), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n694), .A2(new_n855), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n737), .A3(new_n685), .A4(new_n857), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n666), .A2(new_n672), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n616), .A2(new_n304), .A3(new_n655), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n718), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n731), .A2(new_n730), .A3(new_n733), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n701), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n861), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n860), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n860), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n716), .B(new_n713), .C1(new_n368), .C2(new_n617), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n629), .A2(new_n757), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n564), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n569), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n451), .A3(new_n365), .A4(new_n643), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n656), .A3(new_n728), .A4(new_n719), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n659), .A2(new_n514), .A3(new_n665), .A4(new_n739), .ZN(new_n883));
  INV_X1    g697(.A(new_n868), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n737), .A3(new_n739), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n755), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n753), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT52), .B1(new_n866), .B2(new_n869), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n874), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n874), .B2(new_n891), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n746), .B2(new_n752), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n882), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n889), .B1(new_n896), .B2(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n874), .A2(new_n891), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n874), .A2(new_n890), .A3(new_n891), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(KEYINPUT53), .A3(new_n901), .A4(new_n888), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n872), .A2(new_n874), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n837), .B(KEYINPUT120), .C1(new_n849), .C2(new_n851), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n854), .A2(new_n898), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(KEYINPUT54), .B2(new_n897), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n854), .A4(new_n908), .ZN(new_n914));
  INV_X1    g728(.A(G952), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n345), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n814), .B(KEYINPUT49), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n563), .A2(new_n636), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n919), .A2(new_n364), .A3(new_n622), .A4(new_n615), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n686), .A3(new_n920), .A4(new_n693), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n345), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n296), .B1(new_n902), .B2(new_n906), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n409), .A2(new_n418), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n424), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n902), .A2(new_n906), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(KEYINPUT122), .A3(G902), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT122), .B1(new_n931), .B2(G902), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n446), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n934), .B2(new_n936), .ZN(G51));
  XOR2_X1   g751(.A(new_n775), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n903), .B1(new_n902), .B2(new_n906), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n907), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n611), .ZN(new_n945));
  INV_X1    g759(.A(new_n774), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n932), .B2(new_n933), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n923), .B1(new_n945), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n932), .B2(new_n933), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n923), .B1(new_n950), .B2(new_n559), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n552), .B(new_n949), .C1(new_n932), .C2(new_n933), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G60));
  AND2_X1   g767(.A1(new_n631), .A2(new_n632), .ZN(new_n954));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT59), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n943), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n941), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n898), .A2(new_n907), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n954), .B1(new_n960), .B2(new_n956), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n959), .A2(new_n961), .A3(new_n923), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT60), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n902), .B2(new_n906), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n352), .B(KEYINPUT125), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n924), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n965), .B2(new_n653), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n965), .A2(new_n969), .A3(new_n653), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n964), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT53), .B1(new_n875), .B2(new_n888), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n894), .A2(KEYINPUT53), .A3(new_n882), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n892), .A2(new_n893), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n923), .B1(new_n980), .B2(new_n966), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n653), .B(new_n976), .C1(new_n977), .C2(new_n979), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n974), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n972), .A2(new_n973), .ZN(new_n985));
  NAND2_X1  g799(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n975), .A2(new_n987), .ZN(G66));
  NOR3_X1   g802(.A1(new_n568), .A2(new_n422), .A3(new_n345), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n882), .B2(new_n345), .ZN(new_n990));
  INV_X1    g804(.A(G898), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n927), .B1(new_n991), .B2(G953), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n990), .B(new_n992), .Z(G69));
  NAND3_X1  g807(.A1(new_n782), .A2(new_n750), .A3(new_n862), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n755), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n794), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n869), .B1(new_n659), .B2(new_n673), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n784), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT127), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n753), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n1000), .A2(G953), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n236), .A2(new_n261), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(new_n548), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n345), .B1(G227), .B2(G900), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n696), .A2(new_n997), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1010));
  OR3_X1    g824(.A1(new_n677), .A2(new_n738), .A3(new_n878), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n784), .B1(new_n368), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n794), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1009), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1014), .B2(new_n345), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1005), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1006), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  INV_X1    g834(.A(new_n882), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1000), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n923), .B1(new_n1022), .B2(new_n286), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1020), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g838(.A(new_n681), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n265), .B2(new_n278), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1027), .B1(new_n897), .B2(new_n1029), .ZN(G57));
endmodule


