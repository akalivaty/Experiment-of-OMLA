

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583;

  XNOR2_X1 U325 ( .A(n430), .B(KEYINPUT54), .ZN(n431) );
  XNOR2_X1 U326 ( .A(n432), .B(n431), .ZN(n448) );
  XNOR2_X1 U327 ( .A(n415), .B(KEYINPUT64), .ZN(n416) );
  XNOR2_X1 U328 ( .A(n420), .B(n308), .ZN(n309) );
  XNOR2_X1 U329 ( .A(n417), .B(n416), .ZN(n542) );
  XNOR2_X1 U330 ( .A(n310), .B(n309), .ZN(n386) );
  XNOR2_X1 U331 ( .A(KEYINPUT122), .B(n451), .ZN(n563) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XNOR2_X1 U334 ( .A(G106GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n293), .B(KEYINPUT74), .ZN(n339) );
  XNOR2_X1 U336 ( .A(G120GAT), .B(G148GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n294), .B(G57GAT), .ZN(n433) );
  XNOR2_X1 U338 ( .A(n339), .B(n433), .ZN(n301) );
  XNOR2_X1 U339 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n295), .B(KEYINPUT73), .ZN(n372) );
  INV_X1 U341 ( .A(n372), .ZN(n299) );
  XOR2_X1 U342 ( .A(KEYINPUT33), .B(KEYINPUT78), .Z(n297) );
  NAND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n302), .B(KEYINPUT31), .Z(n310) );
  XOR2_X1 U348 ( .A(G92GAT), .B(G64GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(G176GAT), .B(n305), .Z(n420) );
  XOR2_X1 U352 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n307) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G85GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n350) );
  XNOR2_X1 U355 ( .A(n350), .B(KEYINPUT32), .ZN(n308) );
  INV_X1 U356 ( .A(KEYINPUT41), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n386), .B(n311), .ZN(n408) );
  XNOR2_X1 U358 ( .A(KEYINPUT107), .B(n408), .ZN(n532) );
  XNOR2_X1 U359 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(KEYINPUT17), .ZN(n313) );
  XOR2_X1 U361 ( .A(n313), .B(KEYINPUT19), .Z(n315) );
  XNOR2_X1 U362 ( .A(G183GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n427) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G176GAT), .Z(n317) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G15GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n427), .B(n318), .ZN(n329) );
  XNOR2_X1 U368 ( .A(G134GAT), .B(G127GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n319), .B(KEYINPUT0), .ZN(n437) );
  XOR2_X1 U370 ( .A(G99GAT), .B(n437), .Z(n321) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(KEYINPUT84), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(n322), .B(KEYINPUT20), .Z(n327) );
  XOR2_X1 U374 ( .A(KEYINPUT86), .B(G71GAT), .Z(n324) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(G113GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n527) );
  XNOR2_X1 U380 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n330), .B(KEYINPUT3), .ZN(n331) );
  XOR2_X1 U382 ( .A(n331), .B(KEYINPUT88), .Z(n333) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(G162GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n445) );
  XOR2_X1 U385 ( .A(G50GAT), .B(G22GAT), .Z(n392) );
  XOR2_X1 U386 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n335) );
  XNOR2_X1 U387 ( .A(KEYINPUT23), .B(G148GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(n392), .B(n336), .Z(n338) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n445), .B(n343), .ZN(n347) );
  XOR2_X1 U396 ( .A(KEYINPUT21), .B(G218GAT), .Z(n345) );
  XNOR2_X1 U397 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(n346), .ZN(n422) );
  XNOR2_X1 U400 ( .A(n347), .B(n422), .ZN(n465) );
  XOR2_X1 U401 ( .A(G29GAT), .B(G43GAT), .Z(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n404) );
  XNOR2_X1 U404 ( .A(n404), .B(n350), .ZN(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U406 ( .A(G50GAT), .B(G134GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n360) );
  XOR2_X1 U409 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n356) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U412 ( .A(G218GAT), .B(G92GAT), .Z(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n362) );
  NAND2_X1 U415 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U417 ( .A(KEYINPUT80), .B(KEYINPUT11), .Z(n364) );
  XNOR2_X1 U418 ( .A(G162GAT), .B(G106GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n554) );
  XNOR2_X1 U421 ( .A(KEYINPUT36), .B(n554), .ZN(n486) );
  XOR2_X1 U422 ( .A(G78GAT), .B(G211GAT), .Z(n368) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G127GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n369), .B(G155GAT), .Z(n371) );
  XOR2_X1 U426 ( .A(G15GAT), .B(KEYINPUT71), .Z(n389) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(n389), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U429 ( .A(n372), .B(KEYINPUT12), .Z(n374) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U432 ( .A(n376), .B(n375), .Z(n384) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G57GAT), .Z(n378) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(G1GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n380) );
  XNOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n578) );
  NOR2_X1 U441 ( .A1(n486), .A2(n578), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT45), .ZN(n387) );
  NAND2_X1 U443 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT113), .ZN(n407) );
  XOR2_X1 U445 ( .A(G197GAT), .B(G141GAT), .Z(n391) );
  XOR2_X1 U446 ( .A(G113GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U447 ( .A(n434), .B(n389), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n398) );
  XOR2_X1 U450 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n395) );
  NAND2_X1 U451 ( .A1(G229GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT68), .B(n396), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U455 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n400) );
  XNOR2_X1 U456 ( .A(KEYINPUT66), .B(KEYINPUT69), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(G36GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n403), .B(G8GAT), .ZN(n424) );
  XNOR2_X1 U461 ( .A(n404), .B(n424), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n573) );
  XNOR2_X1 U463 ( .A(n573), .B(KEYINPUT72), .ZN(n557) );
  NAND2_X1 U464 ( .A1(n407), .A2(n557), .ZN(n414) );
  NAND2_X1 U465 ( .A1(n578), .A2(n554), .ZN(n411) );
  NOR2_X1 U466 ( .A1(n573), .A2(n408), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT46), .ZN(n410) );
  NOR2_X1 U468 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n412), .B(KEYINPUT47), .ZN(n413) );
  NAND2_X1 U470 ( .A1(n414), .A2(n413), .ZN(n417) );
  INV_X1 U471 ( .A(KEYINPUT48), .ZN(n415) );
  XOR2_X1 U472 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n419) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U475 ( .A(n421), .B(n420), .Z(n426) );
  INV_X1 U476 ( .A(n422), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n518) );
  XOR2_X1 U480 ( .A(n518), .B(KEYINPUT119), .Z(n429) );
  NOR2_X1 U481 ( .A1(n542), .A2(n429), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n430) );
  XOR2_X1 U483 ( .A(n433), .B(G85GAT), .Z(n436) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n436), .B(n435), .ZN(n441) );
  XOR2_X1 U486 ( .A(n437), .B(KEYINPUT1), .Z(n439) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U488 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U489 ( .A(n441), .B(n440), .Z(n447) );
  XOR2_X1 U490 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n443) );
  XNOR2_X1 U491 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n442) );
  XNOR2_X1 U492 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U494 ( .A(n447), .B(n446), .ZN(n469) );
  XNOR2_X1 U495 ( .A(KEYINPUT91), .B(n469), .ZN(n541) );
  NAND2_X1 U496 ( .A1(n448), .A2(n541), .ZN(n570) );
  NOR2_X1 U497 ( .A1(n465), .A2(n570), .ZN(n449) );
  XNOR2_X1 U498 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NOR2_X1 U499 ( .A1(n527), .A2(n450), .ZN(n451) );
  NAND2_X1 U500 ( .A1(n532), .A2(n563), .ZN(n455) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U502 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n452) );
  INV_X1 U503 ( .A(n386), .ZN(n456) );
  NOR2_X1 U504 ( .A1(n456), .A2(n557), .ZN(n491) );
  XOR2_X1 U505 ( .A(n518), .B(KEYINPUT27), .Z(n457) );
  XNOR2_X1 U506 ( .A(n457), .B(KEYINPUT94), .ZN(n463) );
  XNOR2_X1 U507 ( .A(KEYINPUT65), .B(KEYINPUT28), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n458), .B(n465), .ZN(n523) );
  NAND2_X1 U509 ( .A1(n463), .A2(n523), .ZN(n459) );
  NOR2_X1 U510 ( .A1(n541), .A2(n459), .ZN(n529) );
  NAND2_X1 U511 ( .A1(n527), .A2(n529), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT95), .ZN(n471) );
  XOR2_X1 U513 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n462) );
  NAND2_X1 U514 ( .A1(n527), .A2(n465), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n571) );
  AND2_X1 U516 ( .A1(n571), .A2(n463), .ZN(n544) );
  NOR2_X1 U517 ( .A1(n527), .A2(n518), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n466), .Z(n467) );
  NOR2_X1 U520 ( .A1(n544), .A2(n467), .ZN(n468) );
  NOR2_X1 U521 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U522 ( .A1(n471), .A2(n470), .ZN(n487) );
  INV_X1 U523 ( .A(n554), .ZN(n564) );
  NOR2_X1 U524 ( .A1(n564), .A2(n578), .ZN(n472) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U526 ( .A1(n487), .A2(n473), .ZN(n474) );
  XOR2_X1 U527 ( .A(KEYINPUT97), .B(n474), .Z(n504) );
  NAND2_X1 U528 ( .A1(n491), .A2(n504), .ZN(n483) );
  NOR2_X1 U529 ( .A1(n541), .A2(n483), .ZN(n475) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n475), .Z(n476) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n518), .A2(n483), .ZN(n478) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U536 ( .A1(n527), .A2(n483), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n523), .A2(n483), .ZN(n485) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1327GAT) );
  NOR2_X1 U543 ( .A1(n486), .A2(n487), .ZN(n488) );
  NAND2_X1 U544 ( .A1(n578), .A2(n488), .ZN(n489) );
  XNOR2_X1 U545 ( .A(KEYINPUT102), .B(n489), .ZN(n490) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n490), .ZN(n515) );
  NAND2_X1 U547 ( .A1(n515), .A2(n491), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n492), .B(KEYINPUT38), .ZN(n501) );
  NOR2_X1 U549 ( .A1(n501), .A2(n541), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U552 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NOR2_X1 U553 ( .A1(n501), .A2(n518), .ZN(n496) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(n496), .Z(n497) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n499) );
  NOR2_X1 U557 ( .A1(n527), .A2(n501), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n501), .A2(n523), .ZN(n502) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(n502), .Z(n503) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  AND2_X1 U563 ( .A1(n573), .A2(n532), .ZN(n516) );
  NAND2_X1 U564 ( .A1(n504), .A2(n516), .ZN(n510) );
  NOR2_X1 U565 ( .A1(n541), .A2(n510), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(n505), .Z(n506) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n518), .A2(n510), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n507), .Z(n508) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n527), .A2(n510), .ZN(n509) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n510), .A2(n523), .ZN(n514) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n512) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n541), .A2(n522), .ZN(n517) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n522), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n542), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n531) );
  NOR2_X1 U592 ( .A1(n557), .A2(n531), .ZN(n530) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  INV_X1 U595 ( .A(n531), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n537), .A2(n532), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  INV_X1 U598 ( .A(n578), .ZN(n561) );
  NAND2_X1 U599 ( .A1(n561), .A2(n537), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n564), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n573), .A2(n553), .ZN(n545) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n553), .A2(n408), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n578), .A2(n553), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(n555), .Z(n556) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT123), .Z(n560) );
  INV_X1 U623 ( .A(n557), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n558), .A2(n563), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n575) );
  INV_X1 U635 ( .A(n570), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n580) );
  NOR2_X1 U637 ( .A1(n573), .A2(n580), .ZN(n574) );
  XOR2_X1 U638 ( .A(n575), .B(n574), .Z(G1352GAT) );
  NOR2_X1 U639 ( .A1(n386), .A2(n580), .ZN(n577) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n486), .A2(n580), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

