//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  OAI221_X1 g044(.A(new_n463), .B1(new_n464), .B2(new_n467), .C1(new_n469), .C2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n461), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n461), .A2(G112), .ZN(new_n480));
  OAI221_X1 g055(.A(new_n477), .B1(new_n478), .B2(new_n467), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT69), .Z(G162));
  NAND2_X1  g057(.A1(new_n474), .A2(new_n475), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G126), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n461), .A2(G114), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n483), .A2(new_n491), .A3(G138), .A4(new_n461), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n468), .A2(new_n494), .A3(G138), .A4(new_n461), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n488), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(KEYINPUT5), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n499), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n498), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n497), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n497), .B2(KEYINPUT71), .ZN(new_n515));
  OR3_X1    g090(.A1(new_n514), .A2(new_n497), .A3(KEYINPUT71), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n502), .A2(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n499), .B1(new_n516), .B2(new_n515), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n509), .A2(new_n524), .A3(G63), .A4(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(G51), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT7), .Z(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n528), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI211_X1 g108(.A(KEYINPUT75), .B(new_n531), .C1(new_n517), .C2(G89), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n526), .B(new_n527), .C1(new_n533), .C2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AND2_X1   g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n509), .B2(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(new_n538), .B2(new_n497), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n517), .A2(G90), .B1(G52), .B2(new_n518), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n502), .B2(new_n508), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n541), .B(G651), .C1(new_n543), .C2(new_n537), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G171));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n518), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n516), .A2(new_n515), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n509), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n509), .A2(G56), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n497), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n517), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n518), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT73), .B1(new_n503), .B2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n507), .B2(G543), .ZN(new_n568));
  AOI211_X1 g143(.A(KEYINPUT73), .B(new_n499), .C1(new_n504), .C2(new_n506), .ZN(new_n569));
  OAI21_X1  g144(.A(G65), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n566), .B1(new_n572), .B2(G651), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n502), .B2(new_n508), .ZN(new_n575));
  INV_X1    g150(.A(new_n571), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n566), .B(G651), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n563), .B(new_n565), .C1(new_n573), .C2(new_n578), .ZN(G299));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n545), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n539), .A2(KEYINPUT79), .A3(new_n540), .A4(new_n544), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G301));
  OAI21_X1  g158(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g161(.A(KEYINPUT80), .B(G651), .C1(new_n509), .C2(G74), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n517), .A2(G87), .B1(G49), .B2(new_n518), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n517), .A2(G86), .B1(G48), .B2(new_n518), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n502), .B2(new_n508), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT81), .Z(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n509), .A2(G60), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n497), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT82), .Z(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n502), .B2(new_n508), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(G92), .B(new_n549), .C1(new_n568), .C2(new_n569), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n518), .A2(G54), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n517), .A2(new_n613), .A3(G92), .ZN(new_n614));
  AND4_X1   g189(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n605), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n605), .B1(G868), .B2(new_n615), .ZN(G321));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT83), .B1(new_n618), .B2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  MUX2_X1   g195(.A(KEYINPUT83), .B(new_n619), .S(new_n620), .Z(G297));
  MUX2_X1   g196(.A(KEYINPUT83), .B(new_n619), .S(new_n620), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OR3_X1    g204(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(new_n467), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(KEYINPUT84), .B1(new_n484), .B2(new_n629), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT15), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2435), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n661), .B(KEYINPUT17), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n661), .B(KEYINPUT86), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n664), .B(new_n669), .C1(new_n666), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT89), .ZN(new_n678));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XOR2_X1   g254(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n682), .A3(new_n676), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  INV_X1    g260(.A(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n675), .A2(new_n676), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n688), .A3(new_n677), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n685), .B(new_n689), .C1(new_n688), .C2(new_n686), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT90), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT90), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  OR3_X1    g270(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n691), .B2(new_n692), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(G229));
  AND2_X1   g276(.A1(KEYINPUT92), .A2(G16), .ZN(new_n702));
  NOR2_X1   g277(.A1(KEYINPUT92), .A2(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n707));
  INV_X1    g282(.A(G20), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n709), .C1(new_n618), .C2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1956), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n710), .ZN(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G4), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n615), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT96), .B(G1348), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n476), .A2(G128), .ZN(new_n722));
  INV_X1    g297(.A(G140), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n461), .A2(G116), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n723), .B2(new_n467), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n705), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n556), .B2(new_n705), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(G1341), .B(new_n734), .C1(new_n556), .C2(new_n705), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND3_X1   g314(.A1(new_n721), .A2(new_n739), .A3(KEYINPUT98), .ZN(new_n740));
  AOI21_X1  g315(.A(KEYINPUT98), .B1(new_n721), .B2(new_n739), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n713), .B(new_n717), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G164), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G27), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2078), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n634), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n476), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT30), .B(G28), .Z(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(G29), .C2(new_n758), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n742), .A2(new_n746), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n634), .A2(G139), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT25), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n763), .C1(new_n461), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  OR2_X1    g342(.A1(new_n637), .A2(new_n728), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n744), .A2(new_n745), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n760), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n705), .A2(G24), .ZN(new_n771));
  XOR2_X1   g346(.A(G290), .B(KEYINPUT93), .Z(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n705), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(G1986), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n728), .A2(G25), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n634), .A2(G131), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT91), .Z(new_n778));
  INV_X1    g353(.A(G119), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n461), .A2(G107), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n484), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(new_n728), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT35), .B(G1991), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT95), .A2(KEYINPUT34), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n710), .A2(G23), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G288), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n796), .A2(G1976), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G1976), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n795), .ZN(new_n800));
  AOI211_X1 g375(.A(KEYINPUT33), .B(new_n793), .C1(G288), .C2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n705), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n705), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1971), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G1971), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n798), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G6), .A2(G16), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n591), .A2(new_n596), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n791), .B(new_n792), .C1(new_n807), .C2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n807), .A2(new_n789), .A3(new_n790), .A4(new_n812), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n788), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(new_n788), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n770), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n710), .A2(G5), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G171), .B2(new_n710), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1961), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT24), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(G34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(G34), .ZN(new_n827));
  AOI21_X1  g402(.A(G29), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n470), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT99), .B(G2084), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G29), .A2(G35), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G162), .B2(G29), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT29), .B(G2090), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n820), .A2(new_n824), .A3(new_n831), .A4(new_n835), .ZN(G150));
  INV_X1    g411(.A(G150), .ZN(G311));
  NAND2_X1  g412(.A1(new_n518), .A2(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n550), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n509), .A2(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n497), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT102), .B(G860), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n553), .A2(new_n554), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G651), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n517), .A2(G81), .B1(new_n518), .B2(new_n547), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n851), .B(new_n852), .C1(new_n843), .C2(new_n840), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n841), .A2(new_n842), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n517), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n855), .B(new_n856), .C1(new_n555), .C2(new_n552), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n611), .A2(new_n609), .A3(new_n614), .A4(new_n612), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n623), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n846), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n849), .B1(new_n866), .B2(new_n867), .ZN(G145));
  XOR2_X1   g443(.A(new_n783), .B(new_n637), .Z(new_n869));
  XNOR2_X1  g444(.A(G164), .B(new_n726), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n765), .B(new_n640), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n869), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G162), .B(new_n470), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n634), .A2(G142), .B1(G130), .B2(new_n476), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n878), .B(new_n879), .C1(G118), .C2(new_n461), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n752), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n874), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n873), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT105), .B(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT106), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n888), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NAND4_X1  g466(.A1(new_n513), .A2(new_n601), .A3(new_n519), .A4(new_n602), .ZN(new_n892));
  INV_X1    g467(.A(new_n519), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n518), .A2(G47), .ZN(new_n894));
  INV_X1    g469(.A(G85), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n550), .B2(new_n895), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n893), .A2(new_n512), .B1(new_n896), .B2(new_n600), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n809), .ZN(new_n899));
  INV_X1    g474(.A(G288), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n897), .A3(G305), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n906));
  NOR2_X1   g481(.A1(G299), .A2(new_n859), .ZN(new_n907));
  INV_X1    g482(.A(new_n563), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n576), .B1(new_n509), .B2(G65), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT78), .B1(new_n909), .B2(new_n497), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n910), .B2(new_n577), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n615), .B1(new_n911), .B2(new_n565), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G299), .A2(new_n859), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n615), .A3(new_n565), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n858), .B(new_n625), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n914), .A2(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT107), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n905), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n905), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n844), .ZN(G331));
  INV_X1    g504(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(G301), .A2(G168), .ZN(new_n931));
  INV_X1    g506(.A(new_n527), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n509), .A2(G89), .A3(new_n549), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT75), .B1(new_n933), .B2(new_n531), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n529), .A2(new_n528), .A3(new_n532), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n545), .B1(new_n936), .B2(new_n526), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n858), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G286), .B1(new_n581), .B2(new_n582), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n853), .A2(new_n857), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n930), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n940), .B2(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n931), .A2(new_n938), .A3(new_n858), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n918), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n946), .A3(new_n904), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n904), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(G37), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n921), .B2(new_n906), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n955));
  INV_X1    g530(.A(new_n906), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT110), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n944), .A3(new_n945), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(new_n930), .C1(new_n939), .C2(new_n942), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n904), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n943), .A2(new_n946), .A3(new_n904), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n964), .A2(new_n885), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT44), .B(new_n951), .C1(new_n966), .C2(new_n950), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT109), .B1(new_n949), .B2(new_n950), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n943), .A2(new_n946), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n963), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n969), .B(KEYINPUT43), .C1(new_n972), .C2(G37), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n964), .A2(new_n950), .A3(new_n885), .A4(new_n965), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n967), .B1(new_n978), .B2(new_n979), .ZN(G397));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n470), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n726), .B(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT113), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n752), .B(G1996), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n783), .A2(new_n786), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n726), .A2(G2067), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n986), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n988), .B2(new_n752), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(KEYINPUT46), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n986), .B2(G1996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  INV_X1    g577(.A(new_n786), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n990), .B1(new_n1003), .B2(new_n784), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(new_n991), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n995), .ZN(new_n1006));
  OR2_X1    g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(new_n986), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT48), .Z(new_n1009));
  AOI211_X1 g584(.A(new_n994), .B(new_n1002), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n493), .A2(new_n495), .ZN(new_n1011));
  INV_X1    g586(.A(new_n488), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n982), .A3(new_n985), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n716), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1018), .A3(new_n1014), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1020));
  INV_X1    g595(.A(G2084), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n985), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(G168), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT126), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G286), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1024), .A2(new_n1032), .A3(new_n1025), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT62), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n591), .B2(new_n596), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT49), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n1037), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1038), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NOR4_X1   g618(.A1(G164), .A2(new_n470), .A3(new_n984), .A4(G1384), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT116), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n985), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(G8), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1039), .A2(new_n1043), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  AND4_X1   g624(.A1(G1976), .A2(new_n586), .A3(new_n589), .A4(new_n587), .ZN(new_n1050));
  AOI211_X1 g625(.A(KEYINPUT52), .B(new_n1050), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G288), .A2(new_n799), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(G166), .B2(new_n1029), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND4_X1  g633(.A1(G303), .A2(new_n1058), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT114), .B(G1971), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1016), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1019), .A2(new_n1020), .A3(new_n1063), .A4(new_n985), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1029), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT117), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1050), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT52), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1053), .A2(new_n1066), .A3(new_n1069), .A4(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1019), .A2(new_n985), .A3(new_n1020), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(KEYINPUT118), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1063), .B1(new_n1077), .B2(KEYINPUT118), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1062), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1062), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(G8), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1016), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(KEYINPUT53), .A3(new_n745), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1077), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1016), .B2(G2078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G301), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1028), .A2(new_n1096), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1035), .A2(new_n1085), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1094), .B1(new_n1034), .B2(KEYINPUT62), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT127), .A3(new_n1085), .A4(new_n1097), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1049), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1067), .A2(new_n1068), .A3(new_n1052), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1074), .A2(new_n1069), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1066), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n799), .A3(new_n900), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1040), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1107), .A2(new_n1108), .B1(new_n1110), .B2(new_n1070), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1030), .A2(G168), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1076), .B1(new_n1065), .B2(KEYINPUT120), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n1116), .B2(new_n1106), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1076), .A3(new_n1114), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1074), .A2(new_n1069), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1053), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1066), .A2(KEYINPUT63), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1112), .A2(new_n1117), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n1085), .B2(new_n1112), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1111), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1087), .A2(G301), .A3(new_n1091), .A4(new_n1089), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT54), .B1(new_n1094), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1092), .A2(G171), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1127), .A2(KEYINPUT54), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1085), .A2(new_n1131), .A3(new_n1034), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(new_n556), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1015), .A2(new_n982), .A3(new_n997), .A4(new_n985), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(new_n736), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1046), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1134), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1133), .B1(new_n1139), .B2(KEYINPUT124), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n911), .A2(KEYINPUT122), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(G299), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n911), .B(new_n565), .C1(KEYINPUT122), .C2(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT56), .B(G2072), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1086), .A2(new_n1149), .B1(new_n1077), .B2(new_n712), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT61), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT125), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1142), .A2(new_n1156), .A3(new_n1153), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1077), .A2(new_n720), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(G2067), .B2(new_n1046), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(new_n859), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1162), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(KEYINPUT60), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1158), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1151), .A2(new_n859), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1152), .B1(new_n1169), .B2(new_n1162), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1132), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1103), .A2(new_n1126), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1005), .B1(G1986), .B2(G290), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n986), .B1(new_n1173), .B2(new_n1007), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1010), .B1(new_n1172), .B2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g750(.A(G227), .B(G229), .C1(new_n887), .C2(new_n889), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n1177), .A2(G319), .A3(new_n656), .A4(new_n975), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


