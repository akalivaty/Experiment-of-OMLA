//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n466), .B2(new_n468), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n467), .B2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n468), .C1(new_n464), .C2(new_n465), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(new_n468), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT71), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT71), .A2(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT6), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n508), .A2(G88), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n507), .B2(new_n504), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n508), .A2(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n515), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n499), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n521), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n508), .A2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n516), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n502), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n513), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n508), .A2(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n502), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n554));
  OR2_X1    g129(.A1(KEYINPUT71), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(KEYINPUT71), .A2(G651), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(G543), .B1(new_n557), .B2(new_n503), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g137(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n561), .B1(new_n516), .B2(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n553), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n516), .B(G53), .C1(new_n560), .C2(new_n561), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n558), .A2(new_n559), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n566), .B(KEYINPUT73), .C1(new_n567), .C2(new_n561), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n527), .B1(new_n557), .B2(new_n503), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G651), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n565), .A2(new_n568), .A3(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n508), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n516), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  OAI211_X1 g154(.A(G86), .B(new_n527), .C1(new_n557), .C2(new_n503), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n526), .B2(new_n499), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n513), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n580), .B(new_n585), .C1(new_n558), .C2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n508), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n516), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n512), .C2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n569), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n502), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(G54), .A2(new_n516), .B1(new_n602), .B2(G651), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n594), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n599), .A2(new_n594), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n593), .B1(new_n607), .B2(new_n592), .ZN(G284));
  AOI21_X1  g183(.A(new_n593), .B1(new_n607), .B2(new_n592), .ZN(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n592), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n592), .B2(G168), .ZN(G297));
  XOR2_X1   g186(.A(G297), .B(KEYINPUT75), .Z(G280));
  XOR2_X1   g187(.A(KEYINPUT76), .B(G559), .Z(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(G860), .B2(new_n613), .ZN(G148));
  NAND2_X1  g189(.A1(new_n546), .A2(new_n592), .ZN(new_n615));
  INV_X1    g190(.A(new_n613), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n605), .B2(new_n606), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n617), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n467), .A2(G135), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT77), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n480), .A2(G123), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n623), .A2(KEYINPUT78), .B1(new_n624), .B2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(KEYINPUT78), .B2(new_n623), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(new_n469), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  INV_X1    g212(.A(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT80), .ZN(new_n645));
  INV_X1    g220(.A(G1341), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n643), .A2(new_n642), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(new_n641), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n645), .B2(new_n649), .ZN(new_n651));
  OAI21_X1  g226(.A(G1348), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G1341), .ZN(new_n654));
  INV_X1    g229(.A(G1348), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n645), .A2(new_n649), .A3(new_n646), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n652), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n652), .B2(new_n657), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n636), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n652), .A2(new_n657), .ZN(new_n666));
  INV_X1    g241(.A(new_n661), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n668), .A2(KEYINPUT81), .A3(G14), .A4(new_n662), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n691), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n692), .A2(KEYINPUT20), .A3(new_n691), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n693), .B1(new_n691), .B2(new_n689), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  AND2_X1   g281(.A1(new_n469), .A2(G105), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT26), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n707), .B(new_n709), .C1(G141), .C2(new_n467), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n480), .A2(G129), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(KEYINPUT93), .C1(G29), .C2(G32), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(KEYINPUT93), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT92), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n467), .A2(G139), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n477), .A2(G127), .ZN(new_n725));
  NAND2_X1  g300(.A1(G115), .A2(G2104), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n468), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n719), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G2072), .Z(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(KEYINPUT24), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n730), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2084), .ZN(new_n738));
  NOR2_X1   g313(.A1(G27), .A2(G29), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G164), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT97), .B(G2078), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n732), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n730), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n730), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n546), .A2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G19), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(G1341), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT30), .B(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n754), .A2(new_n730), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n628), .B2(new_n730), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n717), .A2(new_n743), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n749), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n749), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n730), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n480), .A2(G128), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(G116), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G2105), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n467), .B2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n773), .A2(KEYINPUT91), .A3(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(KEYINPUT91), .B1(new_n773), .B2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n767), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G5), .A2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT96), .Z(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G301), .B2(new_n749), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n752), .A2(G1341), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n763), .C2(new_n762), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n765), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G4), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n607), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n749), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT98), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n760), .A2(new_n786), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT86), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT87), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n797), .A2(KEYINPUT86), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n797), .A2(KEYINPUT86), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n803), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(G288), .A2(G16), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n749), .A2(G23), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT88), .Z(new_n810));
  AND2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n749), .A2(G22), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G303), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1971), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n802), .A2(new_n805), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G1971), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n815), .A2(new_n820), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(new_n811), .C2(new_n812), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n824), .A2(KEYINPUT89), .A3(new_n805), .A4(new_n802), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n819), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n819), .B2(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n480), .A2(G119), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G107), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n467), .B2(G131), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G29), .ZN(new_n838));
  OR2_X1    g413(.A1(G25), .A2(G29), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT84), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(KEYINPUT84), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT85), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n749), .B1(G290), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(G290), .ZN(new_n849));
  INV_X1    g424(.A(G24), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(G16), .B2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(G1986), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(G1986), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT90), .B1(new_n830), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n817), .A2(new_n818), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT34), .B1(new_n856), .B2(new_n825), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT90), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n829), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT36), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n830), .A2(KEYINPUT90), .A3(new_n854), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n829), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n796), .B1(new_n862), .B2(new_n867), .ZN(G311));
  AOI21_X1  g443(.A(new_n866), .B1(new_n865), .B2(new_n829), .ZN(new_n869));
  AOI211_X1 g444(.A(KEYINPUT36), .B(new_n828), .C1(new_n863), .C2(new_n864), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n795), .B1(new_n869), .B2(new_n870), .ZN(G150));
  NAND2_X1  g446(.A1(new_n508), .A2(G93), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n516), .A2(G55), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n526), .B2(new_n499), .ZN(new_n875));
  AND2_X1   g450(.A1(G80), .A2(G543), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n513), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT99), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n875), .A2(new_n876), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(new_n513), .B1(new_n516), .B2(G55), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n872), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n546), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n546), .A2(new_n878), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n607), .A2(G559), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  AOI21_X1  g469(.A(G860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(G145));
  XNOR2_X1  g475(.A(new_n486), .B(G160), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n627), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n494), .A2(new_n496), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n495), .A4(new_n490), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n497), .A2(KEYINPUT101), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n480), .A2(G130), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n467), .A2(G142), .ZN(new_n909));
  OAI21_X1  g484(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G118), .B2(new_n468), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n908), .B(new_n909), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n632), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n710), .A2(new_n711), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(new_n773), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n773), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n837), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n712), .A2(new_n768), .A3(new_n772), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n773), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n836), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n915), .B1(new_n919), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n907), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n922), .ZN(new_n926));
  INV_X1    g501(.A(new_n915), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n907), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n925), .A2(new_n728), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n728), .B1(new_n925), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n902), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n923), .A2(new_n924), .A3(new_n907), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n729), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n902), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n925), .A2(new_n931), .A3(new_n728), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  XOR2_X1   g519(.A(G303), .B(G288), .Z(new_n945));
  XOR2_X1   g520(.A(G290), .B(G305), .Z(new_n946));
  XOR2_X1   g521(.A(new_n945), .B(new_n946), .Z(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n606), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n613), .B1(new_n949), .B2(new_n604), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n547), .B1(new_n879), .B2(new_n883), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n888), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n599), .A2(new_n603), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n566), .B1(new_n567), .B2(new_n561), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n573), .B1(new_n957), .B2(new_n553), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n958), .A3(new_n568), .ZN(new_n959));
  NAND2_X1  g534(.A1(G299), .A2(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n950), .A2(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n954), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT41), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n956), .B1(new_n958), .B2(new_n568), .ZN(new_n966));
  NOR2_X1   g541(.A1(G299), .A2(new_n955), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT41), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n617), .A2(new_n890), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n965), .B(new_n968), .C1(new_n969), .C2(new_n953), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n963), .B2(new_n970), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n948), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n963), .A2(new_n970), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n947), .A3(new_n972), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G868), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n884), .A2(new_n592), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n944), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n981), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT103), .B(new_n983), .C1(new_n979), .C2(G868), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(G295));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n981), .ZN(G331));
  NAND2_X1  g561(.A1(G301), .A2(KEYINPUT104), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n532), .A2(new_n533), .A3(new_n537), .A4(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(G168), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(G286), .A2(G301), .A3(KEYINPUT104), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n951), .B2(new_n888), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n887), .A2(new_n990), .A3(new_n889), .A4(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n965), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n964), .B1(new_n959), .B2(new_n960), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n995), .B(KEYINPUT105), .C1(new_n996), .C2(new_n997), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n995), .A2(new_n961), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1000), .A2(new_n948), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n935), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n995), .A2(new_n961), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n998), .B2(new_n999), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n948), .B1(new_n1006), .B2(new_n1001), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n996), .A2(KEYINPUT106), .A3(new_n997), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n995), .B1(new_n968), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1002), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n947), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1003), .A3(new_n1015), .A4(new_n935), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1008), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1003), .A3(new_n935), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1014), .A2(new_n1003), .A3(KEYINPUT107), .A4(new_n935), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT43), .A3(new_n1021), .ZN(new_n1022));
  OR3_X1    g597(.A1(new_n1004), .A2(new_n1007), .A3(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1017), .B1(new_n1024), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n497), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT108), .B(G40), .Z(new_n1028));
  NAND3_X1  g603(.A1(new_n470), .A2(new_n474), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G61), .B1(new_n500), .B2(new_n501), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n512), .B1(new_n1031), .B2(new_n583), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(G48), .B2(new_n516), .ZN(new_n1033));
  OAI21_X1  g608(.A(G1981), .B1(new_n1032), .B2(KEYINPUT112), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n580), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n585), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1030), .B1(new_n1040), .B2(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(KEYINPUT49), .C1(new_n1035), .C2(new_n1039), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(G288), .A2(G1976), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(G1981), .B2(G305), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1030), .B(KEYINPUT114), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT109), .B1(new_n1027), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(KEYINPUT45), .C1(new_n497), .C2(new_n1026), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1055), .A2(new_n1057), .A3(new_n1029), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n905), .A2(KEYINPUT45), .A3(new_n906), .A4(new_n1026), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1971), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1029), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n497), .A2(new_n1064), .A3(new_n1026), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT110), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1029), .B1(KEYINPUT50), .B2(new_n1027), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1053), .B1(new_n1060), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1027), .A2(new_n1054), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1056), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1026), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1029), .B1(new_n1078), .B2(KEYINPUT109), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n1059), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n820), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT111), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1072), .A2(G8), .A3(new_n1075), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1027), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1062), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n576), .A2(new_n577), .A3(G1976), .A4(new_n578), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(G8), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1088), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1047), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1052), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1081), .A2(new_n1066), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1096), .B2(new_n1074), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1077), .A2(new_n1079), .A3(new_n1098), .A4(new_n1059), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1068), .A2(new_n1065), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1099), .A2(new_n1100), .B1(new_n782), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1076), .A2(KEYINPUT115), .A3(new_n1062), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1078), .B2(new_n1029), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1084), .A2(KEYINPUT45), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1098), .A2(KEYINPUT53), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G301), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1097), .A2(new_n1083), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  INV_X1    g687(.A(G8), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G168), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1107), .A2(new_n763), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n1113), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1117), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1107), .A2(new_n763), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(G2084), .B2(new_n1101), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1114), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1114), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n1116), .C1(new_n1120), .C2(new_n1113), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1122), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1111), .B1(KEYINPUT62), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1125), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1113), .B(new_n1116), .C1(new_n1120), .C2(G168), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n1130), .A2(KEYINPUT62), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1094), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1097), .A2(new_n1083), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G301), .B(KEYINPUT54), .ZN(new_n1136));
  NAND4_X1  g711(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n1098), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n1026), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(new_n1054), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(new_n1059), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1135), .A2(new_n1136), .B1(new_n1140), .B2(new_n1102), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1134), .A2(KEYINPUT123), .A3(new_n1128), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1097), .A3(new_n1083), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1084), .A2(new_n1062), .A3(new_n777), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1119), .B2(G1348), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n607), .B1(new_n1150), .B2(KEYINPUT60), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1101), .A2(new_n655), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1152), .A2(new_n1149), .B1(new_n605), .B2(new_n606), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1148), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n607), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1155), .B(new_n1147), .C1(new_n1157), .C2(new_n607), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT57), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n563), .A2(new_n564), .B1(new_n573), .B2(KEYINPUT117), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n565), .A2(new_n568), .A3(KEYINPUT57), .A4(new_n574), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1956), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1101), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1077), .A2(new_n1079), .A3(new_n1059), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1165), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT61), .B1(new_n1170), .B2(KEYINPUT120), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1174), .ZN(new_n1177));
  INV_X1    g752(.A(G1996), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1077), .A2(new_n1079), .A3(new_n1178), .A4(new_n1059), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT58), .B(G1341), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1085), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n546), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1182), .B(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1159), .A2(new_n1176), .A3(new_n1177), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1174), .B1(new_n1170), .B2(new_n1153), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1142), .A2(new_n1146), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1097), .A2(new_n1083), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1121), .A2(G168), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR4_X1   g770(.A1(new_n1120), .A2(new_n1192), .A3(new_n1113), .A4(G286), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1083), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1072), .A2(G8), .A3(new_n1082), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1093), .B1(new_n1198), .B2(new_n1074), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1197), .B1(new_n1199), .B2(KEYINPUT116), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT116), .ZN(new_n1201));
  AOI211_X1 g776(.A(new_n1201), .B(new_n1093), .C1(new_n1198), .C2(new_n1074), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1195), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1133), .A2(new_n1191), .A3(new_n1203), .ZN(new_n1204));
  AOI211_X1 g779(.A(KEYINPUT45), .B(new_n1029), .C1(new_n907), .C2(new_n1026), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n916), .B(new_n1178), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n773), .B(new_n777), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n837), .A2(new_n845), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n837), .A2(new_n845), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(G290), .B(G1986), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1205), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1204), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1205), .A2(new_n1178), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT46), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1207), .A2(new_n712), .ZN(new_n1216));
  AOI22_X1  g791(.A1(new_n1214), .A2(new_n1215), .B1(new_n1216), .B2(new_n1205), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1218));
  AND2_X1   g793(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT47), .Z(new_n1222));
  XNOR2_X1  g797(.A(new_n1209), .B(KEYINPUT124), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1224));
  OAI22_X1  g799(.A1(new_n1223), .A2(new_n1224), .B1(G2067), .B2(new_n773), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1205), .ZN(new_n1226));
  NOR2_X1   g801(.A1(G290), .A2(G1986), .ZN(new_n1227));
  AOI21_X1  g802(.A(KEYINPUT48), .B1(new_n1205), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1210), .A2(new_n1205), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1205), .A2(KEYINPUT48), .A3(new_n1227), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1226), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1222), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1213), .A2(new_n1233), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g809(.A1(G227), .A2(new_n462), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n670), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n670), .A2(KEYINPUT126), .A3(new_n1236), .ZN(new_n1240));
  NAND4_X1  g814(.A1(new_n1239), .A2(new_n942), .A3(new_n705), .A4(new_n1240), .ZN(new_n1241));
  AND2_X1   g815(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1242));
  NOR2_X1   g816(.A1(new_n1241), .A2(new_n1242), .ZN(G308));
  OR2_X1    g817(.A1(new_n1241), .A2(new_n1242), .ZN(G225));
endmodule


