//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT96), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(KEYINPUT96), .A3(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  AOI21_X1  g010(.A(G1gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(new_n210), .B2(KEYINPUT97), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n210), .A2(KEYINPUT97), .A3(new_n214), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n215), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(KEYINPUT97), .A3(new_n214), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n212), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  OR2_X1    g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT101), .ZN(new_n226));
  INV_X1    g025(.A(G57gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G64gat), .ZN(new_n228));
  INV_X1    g027(.A(G64gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G57gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n228), .A2(new_n230), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT101), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n233), .A3(new_n224), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(KEYINPUT99), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT99), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G71gat), .A3(G78gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n238), .A3(new_n223), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n232), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n236), .A2(new_n238), .A3(new_n223), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n231), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n229), .A2(G57gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n227), .A2(G64gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT100), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n235), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n221), .B1(new_n222), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n222), .ZN(new_n252));
  NAND2_X1  g051(.A1(G231gat), .A2(G233gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n251), .B(new_n254), .Z(new_n255));
  XOR2_X1   g054(.A(G183gat), .B(G211gat), .Z(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G127gat), .B(G155gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT17), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT14), .ZN(new_n266));
  INV_X1    g065(.A(G29gat), .ZN(new_n267));
  INV_X1    g066(.A(G36gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT93), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(G29gat), .A2(G36gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT94), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G43gat), .B(G50gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT15), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT95), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n279), .A2(KEYINPUT15), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n284), .A2(new_n280), .A3(new_n271), .A4(new_n277), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n282), .B2(new_n285), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n265), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT17), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT104), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G85gat), .A3(G92gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT7), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n293), .A2(new_n296), .A3(G85gat), .A4(G92gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  INV_X1    g098(.A(G85gat), .ZN(new_n300));
  INV_X1    g099(.A(G92gat), .ZN(new_n301));
  AOI22_X1  g100(.A1(KEYINPUT8), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G99gat), .B(G106gat), .Z(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n298), .A3(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT105), .Z(new_n309));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n288), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n286), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n308), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G190gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n310), .B2(new_n316), .ZN(new_n321));
  XNOR2_X1  g120(.A(G134gat), .B(G162gat), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT106), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(KEYINPUT106), .ZN(new_n327));
  OR4_X1    g126(.A1(new_n320), .A2(new_n321), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n320), .B2(new_n321), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n264), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G197gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT11), .B(G169gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT12), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n289), .A2(new_n221), .A3(new_n291), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n220), .A3(new_n217), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n314), .A2(new_n221), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n342), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n339), .B(KEYINPUT13), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n343), .A2(KEYINPUT18), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n343), .A2(KEYINPUT18), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n341), .A2(new_n342), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n339), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT18), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n344), .A2(new_n342), .ZN(new_n354));
  INV_X1    g153(.A(new_n346), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(KEYINPUT18), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n337), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n349), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n349), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G230gat), .A2(G233gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n242), .A2(KEYINPUT100), .A3(new_n246), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n240), .B1(new_n232), .B2(new_n239), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(new_n305), .A3(new_n235), .A4(new_n307), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n248), .A2(new_n308), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n368), .A3(new_n367), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT107), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n367), .A2(KEYINPUT107), .A3(new_n368), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n363), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n370), .A2(new_n367), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n363), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G120gat), .B(G148gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G176gat), .B(G204gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT108), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n380), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(KEYINPUT108), .A3(new_n380), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G64gat), .B(G92gat), .Z(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G197gat), .B(G204gat), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT76), .ZN(new_n399));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G183gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT27), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G183gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT28), .B1(new_n407), .B2(G190gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT66), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n404), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n413), .A3(KEYINPUT67), .ZN(new_n418));
  INV_X1    g217(.A(G169gat), .ZN(new_n419));
  INV_X1    g218(.A(G176gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT68), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(KEYINPUT26), .B2(new_n421), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425));
  INV_X1    g224(.A(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT24), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(new_n417), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT23), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT23), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(G169gat), .B2(G176gat), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n432), .B(new_n434), .C1(new_n419), .C2(new_n420), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n425), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n427), .A2(new_n437), .B1(new_n430), .B2(new_n417), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n437), .B2(new_n427), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n428), .B(KEYINPUT64), .Z(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n435), .A2(new_n425), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n444), .A2(new_n446), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n402), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n424), .A2(new_n443), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT77), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n401), .B(new_n453), .C1(new_n455), .C2(new_n446), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n393), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(KEYINPUT37), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n401), .B1(new_n449), .B2(new_n450), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n402), .B(new_n453), .C1(new_n455), .C2(new_n446), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(KEYINPUT89), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT90), .B(KEYINPUT37), .C1(new_n467), .C2(new_n468), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n459), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n461), .A2(KEYINPUT91), .A3(KEYINPUT38), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n476));
  XNOR2_X1  g275(.A(G113gat), .B(G120gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(KEYINPUT1), .ZN(new_n478));
  XOR2_X1   g277(.A(G127gat), .B(G134gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G155gat), .B(G162gat), .Z(new_n482));
  INV_X1    g281(.A(G148gat), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n483), .A2(KEYINPUT82), .A3(G141gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G141gat), .B(G148gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  INV_X1    g286(.A(G155gat), .ZN(new_n488));
  INV_X1    g287(.A(G162gat), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT2), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n485), .A2(new_n487), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT81), .B(KEYINPUT2), .Z(new_n494));
  OAI21_X1  g293(.A(new_n482), .B1(new_n494), .B2(new_n486), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n481), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G225gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n476), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT84), .B(KEYINPUT3), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n481), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(KEYINPUT3), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n496), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n480), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT4), .B1(new_n481), .B2(new_n496), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n500), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT85), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n515), .A2(new_n476), .A3(new_n506), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(new_n300), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT0), .B(G57gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524));
  INV_X1    g323(.A(new_n522), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n513), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(KEYINPUT6), .A3(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n392), .B1(new_n451), .B2(new_n456), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n464), .A2(new_n474), .A3(new_n475), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G228gat), .A2(G233gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n401), .B1(new_n447), .B2(new_n503), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT29), .B1(new_n398), .B2(new_n400), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n400), .B2(new_n398), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n507), .B1(new_n502), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n533), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n534), .A2(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(KEYINPUT87), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(G228gat), .A3(G233gat), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT86), .B1(new_n401), .B2(new_n447), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT3), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n401), .A2(KEYINPUT86), .A3(new_n447), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n507), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n538), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G78gat), .B(G106gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n203), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G50gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n546), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n504), .A2(new_n505), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n515), .A2(new_n552), .A3(new_n516), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n499), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(KEYINPUT39), .C1(new_n499), .C2(new_n497), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n556), .A3(new_n499), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n525), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n555), .A2(new_n525), .A3(new_n562), .A4(new_n557), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n561), .A2(new_n523), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n530), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n451), .A2(new_n456), .A3(new_n392), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT80), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n451), .A2(new_n569), .A3(new_n456), .A4(new_n392), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n551), .B1(new_n564), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n532), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n457), .A2(new_n393), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n565), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n530), .A2(KEYINPUT30), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n571), .A2(new_n576), .A3(new_n529), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n551), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT69), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n454), .A2(new_n480), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n444), .A2(new_n481), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G227gat), .ZN(new_n584));
  INV_X1    g383(.A(G233gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G99gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(G15gat), .B(G43gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n583), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(KEYINPUT33), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n580), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n583), .B2(new_n586), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n581), .B(new_n582), .C1(new_n584), .C2(new_n585), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n596), .A2(KEYINPUT69), .A3(KEYINPUT33), .A4(new_n591), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n597), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n594), .B2(new_n596), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n600), .B1(new_n605), .B2(KEYINPUT73), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT36), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n597), .A2(new_n601), .A3(KEYINPUT74), .A4(new_n603), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n605), .B2(new_n600), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n600), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n579), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n574), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n607), .ZN(new_n618));
  INV_X1    g417(.A(new_n551), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT35), .B1(new_n620), .B2(new_n578), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n578), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n551), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT35), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n566), .A2(KEYINPUT92), .A3(new_n529), .A4(new_n571), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n331), .B(new_n387), .C1(new_n617), .C2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n529), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g432(.A1(new_n630), .A2(new_n572), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT16), .B(G8gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT110), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n634), .A2(KEYINPUT42), .A3(new_n635), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT111), .Z(new_n642));
  OR2_X1    g441(.A1(new_n634), .A2(new_n214), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(G1325gat));
  NAND2_X1  g443(.A1(new_n608), .A2(new_n614), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n202), .B1(new_n630), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n624), .A2(G15gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n630), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT112), .Z(G1326gat));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n551), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n330), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n621), .A2(new_n628), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n615), .B1(new_n532), .B2(new_n573), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(new_n264), .A3(new_n387), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n267), .A3(new_n631), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT45), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT113), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n330), .B1(new_n617), .B2(new_n629), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(KEYINPUT113), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n656), .A2(new_n661), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n349), .A2(new_n358), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n386), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n264), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n529), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n674), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n657), .A2(new_n268), .A3(new_n572), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT46), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT114), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n572), .ZN(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n673), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n679), .B(new_n681), .C1(KEYINPUT46), .C2(new_n676), .ZN(G1329gat));
  NOR2_X1   g481(.A1(new_n624), .A2(G43gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n657), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT115), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n657), .A2(KEYINPUT115), .A3(new_n683), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n645), .ZN(new_n689));
  OAI21_X1  g488(.A(G43gat), .B1(new_n673), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT116), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n688), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g493(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n686), .A2(new_n687), .ZN(new_n696));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n672), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n666), .B2(new_n667), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(new_n645), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n693), .A2(new_n701), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n657), .B2(new_n551), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n551), .A2(G50gat), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g505(.A1(new_n617), .A2(new_n629), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n331), .A2(new_n669), .A3(new_n386), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n529), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n227), .ZN(G1332gat));
  XNOR2_X1  g510(.A(new_n572), .B(KEYINPUT117), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(G1333gat));
  NOR3_X1   g516(.A1(new_n709), .A2(G71gat), .A3(new_n624), .ZN(new_n718));
  INV_X1    g517(.A(new_n709), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n645), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(G71gat), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n551), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n264), .A2(new_n669), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n386), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n668), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n300), .A3(new_n529), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n656), .B2(KEYINPUT118), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT118), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n663), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT119), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n725), .B1(new_n663), .B2(new_n731), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n656), .A2(KEYINPUT118), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n733), .A3(KEYINPUT119), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n734), .A2(new_n739), .A3(new_n631), .A4(new_n671), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n729), .B1(new_n740), .B2(new_n300), .ZN(G1336gat));
  NOR2_X1   g540(.A1(new_n712), .A2(G92gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n734), .A2(new_n739), .A3(new_n671), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G92gat), .B1(new_n728), .B2(new_n712), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n386), .B(new_n726), .C1(new_n666), .C2(new_n667), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n301), .B1(new_n747), .B2(new_n572), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n671), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n738), .B2(new_n733), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT52), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(G1337gat));
  NOR2_X1   g551(.A1(new_n624), .A2(G99gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n734), .A2(new_n739), .A3(new_n671), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G99gat), .B1(new_n728), .B2(new_n689), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1338gat));
  XOR2_X1   g555(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n757));
  AOI21_X1  g556(.A(new_n661), .B1(new_n656), .B2(new_n664), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n663), .A2(new_n662), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n551), .B(new_n727), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n760), .B2(G106gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n734), .A2(new_n739), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n619), .A2(new_n386), .A3(G106gat), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT121), .Z(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n760), .A2(KEYINPUT120), .A3(G106gat), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT120), .B1(new_n760), .B2(G106gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n738), .B2(new_n733), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n264), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n375), .A2(KEYINPUT54), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n373), .A2(new_n374), .A3(new_n363), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT123), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n373), .A2(new_n363), .A3(new_n374), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n375), .A3(new_n777), .A4(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n380), .B1(new_n375), .B2(KEYINPUT54), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT55), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n783), .B(new_n780), .C1(new_n775), .C2(new_n778), .ZN(new_n784));
  INV_X1    g583(.A(new_n381), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n669), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n354), .A2(new_n355), .B1(new_n350), .B2(new_n339), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n336), .ZN(new_n789));
  AND4_X1   g588(.A1(new_n358), .A2(new_n384), .A3(new_n385), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n653), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n358), .A2(new_n789), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n786), .A2(new_n653), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n772), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n264), .A2(new_n330), .A3(new_n670), .A4(new_n386), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n625), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n631), .A3(new_n712), .ZN(new_n799));
  INV_X1    g598(.A(new_n362), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n529), .B1(new_n795), .B2(new_n796), .ZN(new_n802));
  INV_X1    g601(.A(new_n620), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n712), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(G113gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n669), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n801), .A2(new_n808), .ZN(G1340gat));
  OAI21_X1  g608(.A(G120gat), .B1(new_n799), .B2(new_n386), .ZN(new_n810));
  INV_X1    g609(.A(G120gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n811), .A3(new_n671), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1341gat));
  INV_X1    g612(.A(G127gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n814), .A3(new_n772), .ZN(new_n815));
  AOI21_X1  g614(.A(G127gat), .B1(new_n806), .B2(new_n264), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1342gat));
  OR4_X1    g616(.A1(G134gat), .A2(new_n804), .A3(new_n572), .A4(new_n330), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n819));
  OAI21_X1  g618(.A(G134gat), .B1(new_n799), .B2(new_n330), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(G1343gat));
  NOR3_X1   g621(.A1(new_n805), .A2(new_n529), .A3(new_n645), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n797), .B2(new_n551), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  INV_X1    g624(.A(new_n361), .ZN(new_n826));
  INV_X1    g625(.A(new_n782), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n780), .B1(new_n775), .B2(new_n778), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n785), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n349), .A2(new_n358), .A3(new_n359), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n653), .B1(new_n831), .B2(new_n791), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n772), .B1(new_n832), .B2(new_n794), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n825), .B(new_n619), .C1(new_n833), .C2(new_n796), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n823), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G141gat), .B1(new_n835), .B2(new_n800), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n645), .A2(new_n619), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n802), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n805), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n800), .A2(G141gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n835), .A2(new_n670), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n843), .A2(G141gat), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(G1344gat));
  XOR2_X1   g645(.A(new_n823), .B(KEYINPUT124), .Z(new_n847));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n331), .A2(new_n362), .A3(new_n671), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n786), .A2(new_n653), .A3(new_n793), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n790), .B1(new_n786), .B2(new_n362), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n653), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n852), .B2(new_n772), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n551), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n849), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n833), .A2(new_n856), .A3(new_n854), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n848), .B(new_n825), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n797), .A2(KEYINPUT57), .A3(new_n551), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n833), .A2(new_n856), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT125), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n853), .A2(new_n854), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n551), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n848), .B1(new_n864), .B2(new_n825), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n671), .B(new_n847), .C1(new_n860), .C2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(G148gat), .B1(new_n835), .B2(new_n386), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n386), .A2(G148gat), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n868), .A2(new_n869), .B1(new_n839), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(G1345gat));
  OR3_X1    g671(.A1(new_n835), .A2(new_n488), .A3(new_n772), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(G155gat), .B1(new_n839), .B2(new_n264), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n835), .B2(new_n330), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n680), .A2(new_n489), .A3(new_n653), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n838), .B2(new_n878), .ZN(G1347gat));
  NOR2_X1   g678(.A1(new_n680), .A2(new_n631), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n798), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n800), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n631), .B(new_n712), .C1(new_n795), .C2(new_n796), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n803), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n419), .A3(new_n669), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n886), .B2(new_n671), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n386), .A2(new_n420), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n881), .B2(new_n890), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n885), .A2(new_n407), .A3(new_n772), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n264), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(G183gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n426), .A3(new_n653), .ZN(new_n897));
  OAI21_X1  g696(.A(G190gat), .B1(new_n882), .B2(new_n330), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(KEYINPUT61), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(KEYINPUT61), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1351gat));
  AND2_X1   g700(.A1(new_n884), .A2(new_n837), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n333), .A3(new_n669), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n689), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n362), .B(new_n905), .C1(new_n860), .C2(new_n865), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  INV_X1    g709(.A(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n911), .A3(new_n671), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT62), .Z(new_n913));
  INV_X1    g712(.A(new_n865), .ZN(new_n914));
  INV_X1    g713(.A(new_n859), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n619), .B1(new_n861), .B2(KEYINPUT125), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(new_n916), .B2(new_n863), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(new_n848), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n386), .B(new_n904), .C1(new_n914), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n913), .B1(new_n911), .B2(new_n919), .ZN(G1353gat));
  INV_X1    g719(.A(G211gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n921), .A3(new_n264), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n264), .B(new_n905), .C1(new_n860), .C2(new_n865), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n902), .B2(new_n653), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n904), .B1(new_n914), .B2(new_n918), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n653), .A2(G218gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G1355gat));
endmodule


