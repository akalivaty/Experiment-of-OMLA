

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775;

  XNOR2_X1 U378 ( .A(n383), .B(n459), .ZN(n552) );
  XNOR2_X1 U379 ( .A(n539), .B(KEYINPUT64), .ZN(n764) );
  XNOR2_X2 U380 ( .A(n622), .B(n428), .ZN(n661) );
  OR2_X2 U381 ( .A1(n734), .A2(G902), .ZN(n458) );
  NAND2_X1 U382 ( .A1(n581), .A2(n423), .ZN(n377) );
  NOR2_X2 U383 ( .A1(n772), .A2(n580), .ZN(n581) );
  NOR2_X2 U384 ( .A1(n744), .A2(n749), .ZN(n434) );
  NOR2_X2 U385 ( .A1(n733), .A2(n749), .ZN(n435) );
  NOR2_X1 U386 ( .A1(n697), .A2(n376), .ZN(n577) );
  NAND2_X2 U387 ( .A1(n676), .A2(n678), .ZN(n616) );
  XNOR2_X2 U388 ( .A(n614), .B(KEYINPUT109), .ZN(n676) );
  NOR2_X2 U389 ( .A1(n730), .A2(n656), .ZN(n533) );
  XNOR2_X2 U390 ( .A(n571), .B(KEYINPUT104), .ZN(n771) );
  NOR2_X2 U391 ( .A1(n570), .A2(n573), .ZN(n571) );
  XNOR2_X2 U392 ( .A(n521), .B(n490), .ZN(n383) );
  XNOR2_X2 U393 ( .A(n518), .B(n517), .ZN(n381) );
  XNOR2_X2 U394 ( .A(KEYINPUT71), .B(G110), .ZN(n517) );
  XNOR2_X2 U395 ( .A(n502), .B(n487), .ZN(n521) );
  NAND2_X1 U396 ( .A1(n460), .A2(n366), .ZN(n655) );
  NOR2_X1 U397 ( .A1(n633), .A2(n632), .ZN(n716) );
  XNOR2_X1 U398 ( .A(n461), .B(KEYINPUT103), .ZN(n635) );
  NAND2_X1 U399 ( .A1(n477), .A2(n481), .ZN(n479) );
  XNOR2_X1 U400 ( .A(n554), .B(G472), .ZN(n663) );
  NOR2_X1 U401 ( .A1(n582), .A2(n584), .ZN(n678) );
  NAND2_X1 U402 ( .A1(n494), .A2(n493), .ZN(n518) );
  INV_X2 U403 ( .A(G143), .ZN(n486) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(G902), .ZN(n543) );
  XNOR2_X2 U405 ( .A(n456), .B(n579), .ZN(n772) );
  XNOR2_X1 U406 ( .A(n635), .B(n432), .ZN(n643) );
  INV_X1 U407 ( .A(KEYINPUT82), .ZN(n432) );
  INV_X1 U408 ( .A(KEYINPUT19), .ZN(n484) );
  AND2_X1 U409 ( .A1(n665), .A2(n403), .ZN(n628) );
  NOR2_X1 U410 ( .A1(n666), .A2(n404), .ZN(n403) );
  INV_X1 U411 ( .A(n617), .ZN(n404) );
  INV_X1 U412 ( .A(KEYINPUT41), .ZN(n615) );
  XNOR2_X1 U413 ( .A(n641), .B(KEYINPUT81), .ZN(n439) );
  AND2_X1 U414 ( .A1(n716), .A2(n402), .ZN(n642) );
  NAND2_X1 U415 ( .A1(n389), .A2(n643), .ZN(n596) );
  OR2_X1 U416 ( .A1(n705), .A2(n721), .ZN(n389) );
  NOR2_X1 U417 ( .A1(n665), .A2(n446), .ZN(n445) );
  OR2_X1 U418 ( .A1(n575), .A2(n604), .ZN(n446) );
  XNOR2_X1 U419 ( .A(n589), .B(KEYINPUT105), .ZN(n451) );
  NAND2_X1 U420 ( .A1(n478), .A2(n479), .ZN(n411) );
  AND2_X1 U421 ( .A1(n483), .A2(n368), .ZN(n478) );
  NAND2_X1 U422 ( .A1(n468), .A2(KEYINPUT2), .ZN(n467) );
  INV_X1 U423 ( .A(n655), .ZN(n468) );
  AND2_X1 U424 ( .A1(n719), .A2(n363), .ZN(n627) );
  XNOR2_X1 U425 ( .A(n516), .B(n515), .ZN(n584) );
  NOR2_X1 U426 ( .A1(G902), .A2(n741), .ZN(n516) );
  NOR2_X1 U427 ( .A1(n773), .A2(n775), .ZN(n397) );
  INV_X1 U428 ( .A(KEYINPUT4), .ZN(n487) );
  INV_X1 U429 ( .A(n635), .ZN(n675) );
  NAND2_X1 U430 ( .A1(n378), .A2(n392), .ZN(n391) );
  INV_X1 U431 ( .A(KEYINPUT44), .ZN(n392) );
  NOR2_X1 U432 ( .A1(n415), .A2(n597), .ZN(n414) );
  NAND2_X1 U433 ( .A1(n412), .A2(n597), .ZN(n419) );
  INV_X1 U434 ( .A(n521), .ZN(n472) );
  XNOR2_X1 U435 ( .A(KEYINPUT77), .B(KEYINPUT91), .ZN(n522) );
  XOR2_X1 U436 ( .A(KEYINPUT90), .B(KEYINPUT18), .Z(n523) );
  XNOR2_X1 U437 ( .A(n395), .B(n645), .ZN(n460) );
  INV_X1 U438 ( .A(n726), .ZN(n650) );
  INV_X1 U439 ( .A(KEYINPUT1), .ZN(n428) );
  INV_X1 U440 ( .A(n583), .ZN(n582) );
  XNOR2_X1 U441 ( .A(n529), .B(n469), .ZN(n756) );
  XNOR2_X1 U442 ( .A(n531), .B(n530), .ZN(n469) );
  XOR2_X1 U443 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n530) );
  XNOR2_X1 U444 ( .A(n564), .B(n562), .ZN(n449) );
  XNOR2_X1 U445 ( .A(G128), .B(G110), .ZN(n564) );
  XNOR2_X1 U446 ( .A(G137), .B(G119), .ZN(n562) );
  XNOR2_X1 U447 ( .A(n504), .B(n431), .ZN(n565) );
  INV_X1 U448 ( .A(KEYINPUT8), .ZN(n431) );
  NOR2_X1 U449 ( .A1(n625), .A2(n484), .ZN(n481) );
  NOR2_X1 U450 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U451 ( .A(n409), .B(n408), .ZN(n572) );
  INV_X1 U452 ( .A(KEYINPUT22), .ZN(n408) );
  NOR2_X1 U453 ( .A1(n587), .A2(n410), .ZN(n409) );
  NAND2_X1 U454 ( .A1(n678), .A2(n424), .ZN(n410) );
  BUF_X1 U455 ( .A(n663), .Z(n429) );
  OR2_X1 U456 ( .A1(n747), .A2(G902), .ZN(n405) );
  NOR2_X1 U457 ( .A1(n572), .A2(n450), .ZN(n592) );
  XNOR2_X1 U458 ( .A(n464), .B(n463), .ZN(n514) );
  XNOR2_X1 U459 ( .A(n510), .B(n465), .ZN(n464) );
  XNOR2_X1 U460 ( .A(n527), .B(n513), .ZN(n463) );
  AND2_X1 U461 ( .A1(n695), .A2(n372), .ZN(n454) );
  INV_X1 U462 ( .A(KEYINPUT121), .ZN(n452) );
  INV_X1 U463 ( .A(KEYINPUT47), .ZN(n402) );
  INV_X1 U464 ( .A(KEYINPUT67), .ZN(n492) );
  OR2_X1 U465 ( .A1(n722), .A2(n462), .ZN(n461) );
  INV_X1 U466 ( .A(n596), .ZN(n415) );
  INV_X1 U467 ( .A(KEYINPUT48), .ZN(n645) );
  OR2_X1 U468 ( .A1(G237), .A2(G902), .ZN(n534) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n498) );
  XNOR2_X1 U470 ( .A(G116), .B(G113), .ZN(n497) );
  XOR2_X1 U471 ( .A(KEYINPUT3), .B(G119), .Z(n531) );
  NOR2_X1 U472 ( .A1(G953), .A2(G237), .ZN(n512) );
  XNOR2_X1 U473 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U474 ( .A(G140), .ZN(n547) );
  XNOR2_X1 U475 ( .A(G107), .B(G104), .ZN(n548) );
  INV_X1 U476 ( .A(G146), .ZN(n459) );
  INV_X1 U477 ( .A(KEYINPUT74), .ZN(n400) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n536) );
  INV_X1 U479 ( .A(KEYINPUT76), .ZN(n442) );
  INV_X1 U480 ( .A(n575), .ZN(n424) );
  INV_X1 U481 ( .A(G953), .ZN(n539) );
  XOR2_X1 U482 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n505) );
  XNOR2_X1 U483 ( .A(G134), .B(G122), .ZN(n387) );
  XNOR2_X1 U484 ( .A(n503), .B(n528), .ZN(n388) );
  XNOR2_X1 U485 ( .A(n511), .B(KEYINPUT98), .ZN(n465) );
  XNOR2_X1 U486 ( .A(G143), .B(G131), .ZN(n511) );
  XNOR2_X1 U487 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U488 ( .A(n422), .B(n371), .ZN(n697) );
  INV_X1 U489 ( .A(KEYINPUT2), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n506), .B(G478), .ZN(n583) );
  XNOR2_X1 U491 ( .A(n566), .B(n447), .ZN(n747) );
  XNOR2_X1 U492 ( .A(n563), .B(n449), .ZN(n448) );
  XNOR2_X1 U493 ( .A(n385), .B(n384), .ZN(n701) );
  NAND2_X1 U494 ( .A1(n565), .A2(G217), .ZN(n384) );
  XNOR2_X1 U495 ( .A(n388), .B(n386), .ZN(n385) );
  XNOR2_X1 U496 ( .A(n505), .B(n387), .ZN(n386) );
  NOR2_X1 U497 ( .A1(n696), .A2(n633), .ZN(n623) );
  NOR2_X1 U498 ( .A1(n433), .A2(n646), .ZN(n630) );
  XNOR2_X1 U499 ( .A(n421), .B(n370), .ZN(n580) );
  AND2_X1 U500 ( .A1(n592), .A2(n574), .ZN(n421) );
  XNOR2_X1 U501 ( .A(n591), .B(KEYINPUT31), .ZN(n721) );
  INV_X1 U502 ( .A(n716), .ZN(n710) );
  XNOR2_X1 U503 ( .A(KEYINPUT107), .B(n624), .ZN(n719) );
  NAND2_X1 U504 ( .A1(n595), .A2(n594), .ZN(n702) );
  XNOR2_X1 U505 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U506 ( .A1(n698), .A2(G953), .ZN(n700) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n698) );
  XNOR2_X1 U508 ( .A(n580), .B(n466), .ZN(G21) );
  INV_X1 U509 ( .A(G119), .ZN(n466) );
  XOR2_X1 U510 ( .A(n551), .B(n550), .Z(n357) );
  AND2_X1 U511 ( .A1(n725), .A2(n634), .ZN(n358) );
  AND2_X1 U512 ( .A1(n644), .A2(n439), .ZN(n359) );
  XNOR2_X1 U513 ( .A(KEYINPUT69), .B(G469), .ZN(n360) );
  XOR2_X1 U514 ( .A(G140), .B(KEYINPUT10), .Z(n361) );
  OR2_X1 U515 ( .A1(n625), .A2(n690), .ZN(n362) );
  NOR2_X1 U516 ( .A1(n626), .A2(n362), .ZN(n363) );
  AND2_X1 U517 ( .A1(n359), .A2(n358), .ZN(n364) );
  XOR2_X1 U518 ( .A(n569), .B(n568), .Z(n365) );
  AND2_X1 U519 ( .A1(n728), .A2(n650), .ZN(n366) );
  AND2_X1 U520 ( .A1(n414), .A2(n702), .ZN(n367) );
  NOR2_X1 U521 ( .A1(n542), .A2(n480), .ZN(n368) );
  AND2_X1 U522 ( .A1(n483), .A2(n482), .ZN(n369) );
  XOR2_X1 U523 ( .A(KEYINPUT32), .B(KEYINPUT79), .Z(n370) );
  XOR2_X1 U524 ( .A(n576), .B(KEYINPUT89), .Z(n371) );
  OR2_X1 U525 ( .A1(n697), .A2(n696), .ZN(n372) );
  XOR2_X1 U526 ( .A(n553), .B(KEYINPUT62), .Z(n373) );
  XOR2_X1 U527 ( .A(n701), .B(KEYINPUT124), .Z(n374) );
  NOR2_X1 U528 ( .A1(n764), .A2(G952), .ZN(n749) );
  INV_X1 U529 ( .A(n749), .ZN(n474) );
  XOR2_X1 U530 ( .A(n659), .B(KEYINPUT88), .Z(n375) );
  XNOR2_X1 U531 ( .A(n514), .B(n398), .ZN(n741) );
  XNOR2_X1 U532 ( .A(n448), .B(n398), .ZN(n447) );
  NAND2_X1 U533 ( .A1(n661), .A2(n660), .ZN(n589) );
  BUF_X1 U534 ( .A(n661), .Z(n394) );
  OR2_X1 U535 ( .A1(n621), .A2(n622), .ZN(n633) );
  INV_X1 U536 ( .A(n590), .ZN(n376) );
  XNOR2_X1 U537 ( .A(n411), .B(KEYINPUT0), .ZN(n587) );
  NAND2_X1 U538 ( .A1(n437), .A2(n474), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n438), .B(n373), .ZN(n437) );
  NAND2_X1 U540 ( .A1(n475), .A2(n474), .ZN(n473) );
  XNOR2_X1 U541 ( .A(n476), .B(n374), .ZN(n475) );
  NAND2_X1 U542 ( .A1(n396), .A2(n364), .ZN(n395) );
  XNOR2_X1 U543 ( .A(n397), .B(KEYINPUT46), .ZN(n396) );
  XNOR2_X1 U544 ( .A(n623), .B(KEYINPUT42), .ZN(n773) );
  NAND2_X1 U545 ( .A1(n423), .A2(n581), .ZN(n598) );
  AND2_X1 U546 ( .A1(n423), .A2(n581), .ZN(n378) );
  XNOR2_X1 U547 ( .A(n382), .B(n390), .ZN(n519) );
  BUF_X1 U548 ( .A(n518), .Z(n379) );
  XNOR2_X1 U549 ( .A(n762), .B(n400), .ZN(n399) );
  NOR2_X2 U550 ( .A1(n417), .A2(n418), .ZN(n599) );
  NAND2_X1 U551 ( .A1(n393), .A2(n391), .ZN(n417) );
  NAND2_X1 U552 ( .A1(n420), .A2(n419), .ZN(n418) );
  BUF_X1 U553 ( .A(n730), .Z(n380) );
  NOR2_X1 U554 ( .A1(n653), .A2(n543), .ZN(n401) );
  OR2_X1 U555 ( .A1(n653), .A2(n762), .ZN(n427) );
  NAND2_X1 U556 ( .A1(n413), .A2(n367), .ZN(n393) );
  BUF_X1 U557 ( .A(n608), .Z(n433) );
  XNOR2_X1 U558 ( .A(n608), .B(KEYINPUT38), .ZN(n680) );
  XNOR2_X1 U559 ( .A(n381), .B(n519), .ZN(n520) );
  XNOR2_X1 U560 ( .A(n381), .B(n549), .ZN(n550) );
  XNOR2_X1 U561 ( .A(n361), .B(n382), .ZN(n398) );
  XNOR2_X2 U562 ( .A(G146), .B(G125), .ZN(n382) );
  XNOR2_X1 U563 ( .A(n383), .B(n398), .ZN(n765) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n390) );
  AND2_X2 U565 ( .A1(n693), .A2(n430), .ZN(n745) );
  NAND2_X1 U566 ( .A1(n401), .A2(n399), .ZN(n657) );
  XNOR2_X2 U567 ( .A(n655), .B(n654), .ZN(n762) );
  XNOR2_X2 U568 ( .A(n405), .B(n365), .ZN(n665) );
  NAND2_X1 U569 ( .A1(n406), .A2(n693), .ZN(n743) );
  AND2_X1 U570 ( .A1(n430), .A2(G475), .ZN(n406) );
  NAND2_X1 U571 ( .A1(n407), .A2(n693), .ZN(n732) );
  AND2_X1 U572 ( .A1(n430), .A2(G210), .ZN(n407) );
  NAND2_X1 U573 ( .A1(n745), .A2(G472), .ZN(n438) );
  NAND2_X1 U574 ( .A1(n745), .A2(G478), .ZN(n476) );
  NAND2_X1 U575 ( .A1(n702), .A2(n596), .ZN(n412) );
  NAND2_X1 U576 ( .A1(n598), .A2(KEYINPUT44), .ZN(n413) );
  NAND2_X1 U577 ( .A1(n377), .A2(n416), .ZN(n420) );
  AND2_X1 U578 ( .A1(n597), .A2(KEYINPUT44), .ZN(n416) );
  XNOR2_X2 U579 ( .A(n651), .B(KEYINPUT75), .ZN(n693) );
  NOR2_X1 U580 ( .A1(n583), .A2(n584), .ZN(n585) );
  XNOR2_X2 U581 ( .A(n458), .B(n360), .ZN(n622) );
  XNOR2_X1 U582 ( .A(n552), .B(n357), .ZN(n734) );
  NAND2_X1 U583 ( .A1(n455), .A2(n454), .ZN(n453) );
  XNOR2_X2 U584 ( .A(n533), .B(n532), .ZN(n608) );
  NAND2_X1 U585 ( .A1(n451), .A2(n450), .ZN(n422) );
  INV_X1 U586 ( .A(n771), .ZN(n423) );
  XNOR2_X1 U587 ( .A(n425), .B(KEYINPUT80), .ZN(n694) );
  NAND2_X1 U588 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U589 ( .A(n394), .ZN(n595) );
  INV_X1 U590 ( .A(n626), .ZN(n450) );
  NAND2_X1 U591 ( .A1(n657), .A2(n658), .ZN(n430) );
  XNOR2_X1 U592 ( .A(n434), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U593 ( .A(n435), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U594 ( .A1(n653), .A2(n467), .ZN(n651) );
  XNOR2_X1 U595 ( .A(n436), .B(n375), .ZN(G57) );
  NAND2_X1 U596 ( .A1(n440), .A2(n442), .ZN(n441) );
  NAND2_X1 U597 ( .A1(n445), .A2(n586), .ZN(n440) );
  NAND2_X1 U598 ( .A1(n443), .A2(n441), .ZN(n607) );
  NAND2_X1 U599 ( .A1(n444), .A2(n445), .ZN(n443) );
  AND2_X1 U600 ( .A1(n586), .A2(KEYINPUT76), .ZN(n444) );
  NAND2_X1 U601 ( .A1(n660), .A2(n586), .ZN(n605) );
  NOR2_X1 U602 ( .A1(n665), .A2(n575), .ZN(n660) );
  NAND2_X1 U603 ( .A1(n694), .A2(n693), .ZN(n455) );
  NAND2_X1 U604 ( .A1(n457), .A2(n578), .ZN(n456) );
  XNOR2_X1 U605 ( .A(n577), .B(KEYINPUT34), .ZN(n457) );
  INV_X1 U606 ( .A(n722), .ZN(n711) );
  INV_X1 U607 ( .A(n624), .ZN(n462) );
  XNOR2_X2 U608 ( .A(n599), .B(KEYINPUT45), .ZN(n653) );
  XNOR2_X1 U609 ( .A(n470), .B(n756), .ZN(n730) );
  XNOR2_X1 U610 ( .A(n471), .B(n526), .ZN(n470) );
  XNOR2_X1 U611 ( .A(n520), .B(n472), .ZN(n471) );
  XNOR2_X1 U612 ( .A(n473), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U613 ( .A1(n608), .A2(n484), .ZN(n483) );
  INV_X1 U614 ( .A(n608), .ZN(n477) );
  NAND2_X1 U615 ( .A1(n369), .A2(n479), .ZN(n632) );
  INV_X1 U616 ( .A(n482), .ZN(n480) );
  NAND2_X1 U617 ( .A1(n625), .A2(n484), .ZN(n482) );
  XNOR2_X1 U618 ( .A(KEYINPUT30), .B(n606), .ZN(n485) );
  XNOR2_X1 U619 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U620 ( .A(n552), .B(n501), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n380), .B(n729), .ZN(n731) );
  XNOR2_X1 U622 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U623 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X2 U624 ( .A(n486), .B(G128), .ZN(n502) );
  XOR2_X1 U625 ( .A(KEYINPUT68), .B(G131), .Z(n489) );
  XNOR2_X1 U626 ( .A(G137), .B(G134), .ZN(n488) );
  XNOR2_X1 U627 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U628 ( .A(G101), .ZN(n491) );
  NAND2_X1 U629 ( .A1(n491), .A2(KEYINPUT67), .ZN(n494) );
  NAND2_X1 U630 ( .A1(n492), .A2(G101), .ZN(n493) );
  XOR2_X1 U631 ( .A(n379), .B(n531), .Z(n496) );
  NAND2_X1 U632 ( .A1(n512), .A2(G210), .ZN(n495) );
  XNOR2_X1 U633 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U634 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U635 ( .A(n502), .B(KEYINPUT7), .ZN(n503) );
  XOR2_X1 U636 ( .A(G116), .B(G107), .Z(n528) );
  NAND2_X1 U637 ( .A1(n764), .A2(G234), .ZN(n504) );
  NOR2_X1 U638 ( .A1(n701), .A2(G902), .ZN(n506) );
  XNOR2_X1 U639 ( .A(G113), .B(G104), .ZN(n507) );
  XNOR2_X1 U640 ( .A(n507), .B(G122), .ZN(n527) );
  XOR2_X1 U641 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n509) );
  XNOR2_X1 U642 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n508) );
  XNOR2_X1 U643 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U644 ( .A1(G214), .A2(n512), .ZN(n513) );
  XNOR2_X1 U645 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  NAND2_X1 U646 ( .A1(G224), .A2(n764), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U648 ( .A(n528), .B(n527), .ZN(n529) );
  INV_X1 U649 ( .A(n543), .ZN(n656) );
  AND2_X1 U650 ( .A1(G210), .A2(n534), .ZN(n532) );
  NAND2_X1 U651 ( .A1(n534), .A2(G214), .ZN(n535) );
  XNOR2_X1 U652 ( .A(KEYINPUT92), .B(n535), .ZN(n679) );
  INV_X1 U653 ( .A(n679), .ZN(n625) );
  XNOR2_X1 U654 ( .A(G898), .B(KEYINPUT93), .ZN(n752) );
  NAND2_X1 U655 ( .A1(G953), .A2(n752), .ZN(n758) );
  XOR2_X1 U656 ( .A(n536), .B(KEYINPUT14), .Z(n690) );
  INV_X1 U657 ( .A(n690), .ZN(n603) );
  NAND2_X1 U658 ( .A1(G902), .A2(n603), .ZN(n537) );
  NOR2_X1 U659 ( .A1(n758), .A2(n537), .ZN(n538) );
  XNOR2_X1 U660 ( .A(n538), .B(KEYINPUT94), .ZN(n541) );
  NAND2_X1 U661 ( .A1(G952), .A2(n539), .ZN(n601) );
  NOR2_X1 U662 ( .A1(n601), .A2(n690), .ZN(n540) );
  NOR2_X1 U663 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U664 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n545) );
  NAND2_X1 U665 ( .A1(G234), .A2(n543), .ZN(n544) );
  XNOR2_X1 U666 ( .A(n545), .B(n544), .ZN(n567) );
  NAND2_X1 U667 ( .A1(n567), .A2(G221), .ZN(n546) );
  XNOR2_X1 U668 ( .A(n546), .B(KEYINPUT21), .ZN(n666) );
  XNOR2_X1 U669 ( .A(n666), .B(KEYINPUT96), .ZN(n575) );
  NAND2_X1 U670 ( .A1(G227), .A2(n764), .ZN(n551) );
  NOR2_X1 U671 ( .A1(n553), .A2(G902), .ZN(n554) );
  NAND2_X1 U672 ( .A1(n595), .A2(n429), .ZN(n555) );
  NOR2_X1 U673 ( .A1(n572), .A2(n555), .ZN(n556) );
  XNOR2_X1 U674 ( .A(n556), .B(KEYINPUT65), .ZN(n570) );
  INV_X1 U675 ( .A(KEYINPUT70), .ZN(n557) );
  NAND2_X1 U676 ( .A1(KEYINPUT24), .A2(n557), .ZN(n560) );
  INV_X1 U677 ( .A(KEYINPUT24), .ZN(n558) );
  NAND2_X1 U678 ( .A1(n558), .A2(KEYINPUT70), .ZN(n559) );
  NAND2_X1 U679 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U680 ( .A(n561), .B(KEYINPUT23), .ZN(n563) );
  NAND2_X1 U681 ( .A1(G221), .A2(n565), .ZN(n566) );
  NAND2_X1 U682 ( .A1(n567), .A2(G217), .ZN(n569) );
  INV_X1 U683 ( .A(KEYINPUT25), .ZN(n568) );
  INV_X1 U684 ( .A(n665), .ZN(n573) );
  XOR2_X1 U685 ( .A(n663), .B(KEYINPUT6), .Z(n626) );
  NOR2_X1 U686 ( .A1(n573), .A2(n595), .ZN(n574) );
  XNOR2_X1 U687 ( .A(KEYINPUT35), .B(KEYINPUT84), .ZN(n579) );
  XOR2_X1 U688 ( .A(KEYINPUT33), .B(KEYINPUT106), .Z(n576) );
  AND2_X1 U689 ( .A1(n582), .A2(n584), .ZN(n638) );
  XNOR2_X1 U690 ( .A(n638), .B(KEYINPUT78), .ZN(n578) );
  NAND2_X1 U691 ( .A1(n584), .A2(n583), .ZN(n624) );
  XNOR2_X1 U692 ( .A(KEYINPUT102), .B(n585), .ZN(n722) );
  INV_X1 U693 ( .A(n622), .ZN(n586) );
  INV_X1 U694 ( .A(n587), .ZN(n590) );
  NAND2_X1 U695 ( .A1(n429), .A2(n590), .ZN(n588) );
  NOR2_X1 U696 ( .A1(n605), .A2(n588), .ZN(n705) );
  NOR2_X1 U697 ( .A1(n429), .A2(n589), .ZN(n672) );
  NAND2_X1 U698 ( .A1(n590), .A2(n672), .ZN(n591) );
  XOR2_X1 U699 ( .A(n592), .B(KEYINPUT86), .Z(n593) );
  NOR2_X1 U700 ( .A1(n665), .A2(n593), .ZN(n594) );
  INV_X1 U701 ( .A(KEYINPUT87), .ZN(n597) );
  NOR2_X1 U702 ( .A1(n764), .A2(G900), .ZN(n600) );
  NAND2_X1 U703 ( .A1(G902), .A2(n600), .ZN(n602) );
  NAND2_X1 U704 ( .A1(n602), .A2(n601), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n603), .A2(n617), .ZN(n604) );
  NOR2_X1 U706 ( .A1(n663), .A2(n625), .ZN(n606) );
  NAND2_X1 U707 ( .A1(n607), .A2(n485), .ZN(n636) );
  INV_X1 U708 ( .A(n636), .ZN(n609) );
  NAND2_X1 U709 ( .A1(n609), .A2(n680), .ZN(n612) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(KEYINPUT72), .ZN(n610) );
  XNOR2_X1 U711 ( .A(n610), .B(KEYINPUT39), .ZN(n611) );
  XNOR2_X1 U712 ( .A(n612), .B(n611), .ZN(n649) );
  NOR2_X1 U713 ( .A1(n649), .A2(n624), .ZN(n613) );
  XNOR2_X1 U714 ( .A(KEYINPUT40), .B(n613), .ZN(n775) );
  NAND2_X1 U715 ( .A1(n679), .A2(n680), .ZN(n614) );
  XNOR2_X2 U716 ( .A(n616), .B(n615), .ZN(n696) );
  INV_X1 U717 ( .A(n628), .ZN(n619) );
  OR2_X1 U718 ( .A1(n663), .A2(n690), .ZN(n618) );
  XOR2_X1 U719 ( .A(KEYINPUT28), .B(n620), .Z(n621) );
  NAND2_X1 U720 ( .A1(n628), .A2(n627), .ZN(n646) );
  XNOR2_X1 U721 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n629) );
  XNOR2_X1 U722 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U723 ( .A1(n394), .A2(n631), .ZN(n725) );
  NAND2_X1 U724 ( .A1(KEYINPUT47), .A2(n710), .ZN(n634) );
  NAND2_X1 U725 ( .A1(n635), .A2(KEYINPUT47), .ZN(n640) );
  NOR2_X1 U726 ( .A1(n433), .A2(n636), .ZN(n637) );
  XNOR2_X1 U727 ( .A(KEYINPUT108), .B(n637), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n715) );
  NAND2_X1 U729 ( .A1(n640), .A2(n715), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n644) );
  OR2_X1 U731 ( .A1(n394), .A2(n646), .ZN(n647) );
  XNOR2_X1 U732 ( .A(n647), .B(KEYINPUT43), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n648), .A2(n433), .ZN(n728) );
  NOR2_X1 U734 ( .A1(n649), .A2(n711), .ZN(n726) );
  NAND2_X1 U735 ( .A1(KEYINPUT2), .A2(n656), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n652), .B(KEYINPUT66), .ZN(n658) );
  INV_X1 U737 ( .A(KEYINPUT83), .ZN(n654) );
  XNOR2_X1 U738 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n659) );
  OR2_X1 U739 ( .A1(n394), .A2(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(KEYINPUT50), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n664), .A2(n429), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n667), .ZN(n668) );
  NOR2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT51), .B(n673), .Z(n674) );
  NOR2_X1 U748 ( .A1(n696), .A2(n674), .ZN(n687) );
  NAND2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U750 ( .A(KEYINPUT119), .B(n677), .ZN(n684) );
  INV_X1 U751 ( .A(n678), .ZN(n682) );
  NOR2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n697), .A2(n685), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  NOR2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U759 ( .A1(G952), .A2(n691), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT120), .ZN(n695) );
  XNOR2_X1 U761 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n700), .B(n699), .ZN(G75) );
  XNOR2_X1 U763 ( .A(G101), .B(KEYINPUT112), .ZN(n703) );
  XNOR2_X1 U764 ( .A(n703), .B(n702), .ZN(G3) );
  NAND2_X1 U765 ( .A1(n705), .A2(n719), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n704), .B(G104), .ZN(G6) );
  XOR2_X1 U767 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n707) );
  NAND2_X1 U768 ( .A1(n705), .A2(n722), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n707), .B(n706), .ZN(n709) );
  XOR2_X1 U770 ( .A(G107), .B(KEYINPUT113), .Z(n708) );
  XNOR2_X1 U771 ( .A(n709), .B(n708), .ZN(G9) );
  NOR2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n713) );
  XNOR2_X1 U773 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n712) );
  XNOR2_X1 U774 ( .A(n713), .B(n712), .ZN(n714) );
  XOR2_X1 U775 ( .A(G128), .B(n714), .Z(G30) );
  XNOR2_X1 U776 ( .A(n715), .B(G143), .ZN(G45) );
  NAND2_X1 U777 ( .A1(n716), .A2(n719), .ZN(n717) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT116), .ZN(n718) );
  XNOR2_X1 U779 ( .A(G146), .B(n718), .ZN(G48) );
  NAND2_X1 U780 ( .A1(n721), .A2(n719), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n720), .B(G113), .ZN(G15) );
  NAND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(n723), .B(G116), .ZN(G18) );
  XOR2_X1 U784 ( .A(G125), .B(KEYINPUT37), .Z(n724) );
  XNOR2_X1 U785 ( .A(n725), .B(n724), .ZN(G27) );
  XNOR2_X1 U786 ( .A(G134), .B(n726), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n727), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U788 ( .A(G140), .B(n728), .ZN(G42) );
  XOR2_X1 U789 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n729) );
  XNOR2_X1 U790 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n734), .B(KEYINPUT57), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n745), .A2(G469), .ZN(n737) );
  XNOR2_X1 U794 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n749), .A2(n739), .ZN(G54) );
  INV_X1 U796 ( .A(KEYINPUT59), .ZN(n740) );
  NAND2_X1 U797 ( .A1(G217), .A2(n745), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U799 ( .A1(n749), .A2(n748), .ZN(G66) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n750) );
  XOR2_X1 U801 ( .A(KEYINPUT61), .B(n750), .Z(n751) );
  NOR2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U803 ( .A1(G953), .A2(n653), .ZN(n753) );
  NOR2_X1 U804 ( .A1(n754), .A2(n753), .ZN(n761) );
  XOR2_X1 U805 ( .A(G110), .B(KEYINPUT126), .Z(n755) );
  XNOR2_X1 U806 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n757), .B(G101), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G69) );
  XOR2_X1 U810 ( .A(n762), .B(n765), .Z(n763) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(n769) );
  XOR2_X1 U812 ( .A(G227), .B(n765), .Z(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U814 ( .A1(G953), .A2(n767), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U816 ( .A(G110), .B(KEYINPUT114), .Z(n770) );
  XNOR2_X1 U817 ( .A(n771), .B(n770), .ZN(G12) );
  XOR2_X1 U818 ( .A(n772), .B(G122), .Z(G24) );
  XNOR2_X1 U819 ( .A(G137), .B(KEYINPUT127), .ZN(n774) );
  XNOR2_X1 U820 ( .A(n774), .B(n773), .ZN(G39) );
  XOR2_X1 U821 ( .A(n775), .B(G131), .Z(G33) );
endmodule

