

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770;

  INV_X1 U370 ( .A(KEYINPUT35), .ZN(n348) );
  XNOR2_X1 U371 ( .A(n414), .B(n418), .ZN(n398) );
  XNOR2_X1 U372 ( .A(n530), .B(n359), .ZN(n686) );
  NOR2_X1 U373 ( .A1(n473), .A2(n692), .ZN(n589) );
  NOR2_X1 U374 ( .A1(n608), .A2(n607), .ZN(n618) );
  XNOR2_X1 U375 ( .A(n521), .B(n472), .ZN(n692) );
  XNOR2_X1 U376 ( .A(n552), .B(n419), .ZN(n527) );
  XNOR2_X1 U377 ( .A(n540), .B(n539), .ZN(n741) );
  XNOR2_X1 U378 ( .A(n476), .B(n475), .ZN(n540) );
  XNOR2_X1 U379 ( .A(n487), .B(n486), .ZN(n553) );
  XNOR2_X1 U380 ( .A(G128), .B(KEYINPUT81), .ZN(n400) );
  NOR2_X1 U381 ( .A1(n347), .A2(n617), .ZN(n465) );
  NAND2_X1 U382 ( .A1(n632), .A2(n495), .ZN(n347) );
  XNOR2_X1 U383 ( .A(n513), .B(n563), .ZN(n644) );
  INV_X2 U384 ( .A(n381), .ZN(n666) );
  XNOR2_X1 U385 ( .A(n533), .B(n496), .ZN(n552) );
  INV_X1 U386 ( .A(n349), .ZN(n766) );
  NAND2_X1 U387 ( .A1(n363), .A2(n349), .ZN(n367) );
  XNOR2_X2 U388 ( .A(n573), .B(n348), .ZN(n349) );
  BUF_X2 U389 ( .A(n473), .Z(n443) );
  NOR2_X1 U390 ( .A1(n671), .A2(n668), .ZN(n708) );
  XNOR2_X1 U391 ( .A(n488), .B(G953), .ZN(n506) );
  XNOR2_X2 U392 ( .A(n634), .B(KEYINPUT38), .ZN(n704) );
  NOR2_X2 U393 ( .A1(n644), .A2(G902), .ZN(n518) );
  NOR2_X1 U394 ( .A1(n692), .A2(n606), .ZN(n601) );
  XNOR2_X2 U395 ( .A(n606), .B(KEYINPUT1), .ZN(n473) );
  INV_X1 U396 ( .A(n616), .ZN(n668) );
  INV_X1 U397 ( .A(n613), .ZN(n576) );
  OR2_X1 U398 ( .A1(n398), .A2(n417), .ZN(n396) );
  AND2_X1 U399 ( .A1(n548), .A2(n597), .ZN(n461) );
  XNOR2_X1 U400 ( .A(n400), .B(G143), .ZN(n533) );
  INV_X1 U401 ( .A(KEYINPUT16), .ZN(n538) );
  INV_X1 U402 ( .A(KEYINPUT64), .ZN(n488) );
  INV_X1 U403 ( .A(G475), .ZN(n375) );
  NOR2_X1 U404 ( .A1(n653), .A2(n739), .ZN(n444) );
  NOR2_X1 U405 ( .A1(n733), .A2(n739), .ZN(n735) );
  XNOR2_X1 U406 ( .A(n470), .B(n469), .ZN(n643) );
  NAND2_X1 U407 ( .A1(n352), .A2(n467), .ZN(n470) );
  OR2_X1 U408 ( .A1(n637), .A2(KEYINPUT87), .ZN(n478) );
  XNOR2_X1 U409 ( .A(n392), .B(n391), .ZN(n390) );
  XNOR2_X1 U410 ( .A(n603), .B(KEYINPUT40), .ZN(n769) );
  NAND2_X1 U411 ( .A1(n454), .A2(n450), .ZN(n767) );
  NOR2_X1 U412 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U413 ( .A1(n416), .A2(KEYINPUT34), .ZN(n415) );
  NOR2_X1 U414 ( .A1(n592), .A2(n591), .ZN(n657) );
  AND2_X1 U415 ( .A1(n600), .A2(n471), .ZN(n625) );
  AND2_X1 U416 ( .A1(n414), .A2(n477), .ZN(n574) );
  NAND2_X1 U417 ( .A1(n589), .A2(n576), .ZN(n530) );
  AND2_X1 U418 ( .A1(n609), .A2(n688), .ZN(n477) );
  XNOR2_X1 U419 ( .A(n598), .B(KEYINPUT6), .ZN(n613) );
  NAND2_X1 U420 ( .A1(n405), .A2(n402), .ZN(n598) );
  XNOR2_X1 U421 ( .A(n413), .B(KEYINPUT72), .ZN(n476) );
  XNOR2_X1 U422 ( .A(n564), .B(n538), .ZN(n539) );
  XNOR2_X1 U423 ( .A(G119), .B(G116), .ZN(n475) );
  INV_X1 U424 ( .A(KEYINPUT71), .ZN(n379) );
  NOR2_X1 U425 ( .A1(n687), .A2(n490), .ZN(n489) );
  NAND2_X1 U426 ( .A1(n688), .A2(n353), .ZN(n490) );
  NOR2_X1 U427 ( .A1(n378), .A2(n613), .ZN(n615) );
  XNOR2_X1 U428 ( .A(n401), .B(n442), .ZN(n459) );
  INV_X1 U429 ( .A(KEYINPUT103), .ZN(n442) );
  OR2_X1 U430 ( .A1(n443), .A2(n687), .ZN(n401) );
  AND2_X1 U431 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U432 ( .A1(G472), .A2(G902), .ZN(n406) );
  XNOR2_X1 U433 ( .A(n432), .B(n491), .ZN(n623) );
  INV_X1 U434 ( .A(n657), .ZN(n428) );
  INV_X1 U435 ( .A(KEYINPUT44), .ZN(n388) );
  NOR2_X1 U436 ( .A1(n582), .A2(n388), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n412), .B(KEYINPUT4), .ZN(n537) );
  INV_X1 U438 ( .A(G146), .ZN(n412) );
  OR2_X1 U439 ( .A1(G237), .A2(G902), .ZN(n546) );
  XNOR2_X1 U440 ( .A(n514), .B(KEYINPUT20), .ZN(n519) );
  XNOR2_X1 U441 ( .A(n537), .B(n385), .ZN(n419) );
  XNOR2_X1 U442 ( .A(n411), .B(G131), .ZN(n385) );
  INV_X1 U443 ( .A(G137), .ZN(n411) );
  XNOR2_X1 U444 ( .A(G140), .B(G104), .ZN(n497) );
  XOR2_X1 U445 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n498) );
  XNOR2_X1 U446 ( .A(n527), .B(n474), .ZN(n753) );
  XNOR2_X1 U447 ( .A(KEYINPUT70), .B(KEYINPUT96), .ZN(n474) );
  XNOR2_X1 U448 ( .A(n500), .B(n522), .ZN(n534) );
  XNOR2_X1 U449 ( .A(n386), .B(n462), .ZN(n637) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n462) );
  INV_X1 U451 ( .A(n770), .ZN(n482) );
  NOR2_X1 U452 ( .A1(n616), .A2(n431), .ZN(n430) );
  INV_X1 U453 ( .A(n703), .ZN(n431) );
  NAND2_X1 U454 ( .A1(G214), .A2(n546), .ZN(n703) );
  INV_X1 U455 ( .A(KEYINPUT69), .ZN(n472) );
  XNOR2_X1 U456 ( .A(n569), .B(n568), .ZN(n730) );
  INV_X1 U457 ( .A(KEYINPUT65), .ZN(n469) );
  NAND2_X1 U458 ( .A1(G237), .A2(G234), .ZN(n531) );
  INV_X1 U459 ( .A(n626), .ZN(n634) );
  OR2_X1 U460 ( .A1(n459), .A2(n576), .ZN(n457) );
  NOR2_X1 U461 ( .A1(n459), .A2(n452), .ZN(n451) );
  XNOR2_X1 U462 ( .A(n426), .B(KEYINPUT99), .ZN(n697) );
  NAND2_X1 U463 ( .A1(n589), .A2(n598), .ZN(n426) );
  BUF_X1 U464 ( .A(n506), .Z(n441) );
  NAND2_X1 U465 ( .A1(n409), .A2(n425), .ZN(n440) );
  INV_X1 U466 ( .A(n443), .ZN(n425) );
  XNOR2_X1 U467 ( .A(n410), .B(n358), .ZN(n409) );
  INV_X1 U468 ( .A(KEYINPUT74), .ZN(n491) );
  XNOR2_X1 U469 ( .A(n440), .B(n439), .ZN(n617) );
  INV_X1 U470 ( .A(KEYINPUT90), .ZN(n439) );
  NAND2_X1 U471 ( .A1(n528), .A2(n404), .ZN(n403) );
  INV_X1 U472 ( .A(G902), .ZN(n404) );
  INV_X1 U473 ( .A(KEYINPUT102), .ZN(n391) );
  NAND2_X1 U474 ( .A1(n365), .A2(n349), .ZN(n364) );
  XNOR2_X1 U475 ( .A(G125), .B(KEYINPUT10), .ZN(n505) );
  NOR2_X1 U476 ( .A1(G953), .A2(G237), .ZN(n565) );
  XNOR2_X1 U477 ( .A(G113), .B(G143), .ZN(n560) );
  XOR2_X1 U478 ( .A(KEYINPUT11), .B(G131), .Z(n561) );
  XNOR2_X1 U479 ( .A(G125), .B(KEYINPUT79), .ZN(n541) );
  XOR2_X1 U480 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n542) );
  XNOR2_X1 U481 ( .A(n399), .B(n492), .ZN(n449) );
  XNOR2_X1 U482 ( .A(n533), .B(n536), .ZN(n399) );
  XOR2_X1 U483 ( .A(KEYINPUT78), .B(KEYINPUT93), .Z(n536) );
  XNOR2_X1 U484 ( .A(n545), .B(n493), .ZN(n626) );
  NOR2_X1 U485 ( .A1(n646), .A2(n544), .ZN(n545) );
  XNOR2_X1 U486 ( .A(n377), .B(n520), .ZN(n688) );
  NAND2_X1 U487 ( .A1(n519), .A2(G221), .ZN(n377) );
  XOR2_X1 U488 ( .A(G110), .B(G107), .Z(n740) );
  XNOR2_X1 U489 ( .A(n509), .B(n351), .ZN(n387) );
  XNOR2_X1 U490 ( .A(n380), .B(KEYINPUT24), .ZN(n509) );
  INV_X1 U491 ( .A(KEYINPUT70), .ZN(n380) );
  INV_X1 U492 ( .A(KEYINPUT8), .ZN(n486) );
  INV_X1 U493 ( .A(G134), .ZN(n496) );
  XNOR2_X1 U494 ( .A(G107), .B(G116), .ZN(n549) );
  XNOR2_X1 U495 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U496 ( .A(n494), .B(n499), .ZN(n502) );
  XNOR2_X1 U497 ( .A(n448), .B(n446), .ZN(n646) );
  XNOR2_X1 U498 ( .A(n534), .B(n447), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n741), .B(n449), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n543), .B(n535), .ZN(n447) );
  NOR2_X1 U501 ( .A1(n483), .A2(n482), .ZN(n481) );
  INV_X1 U502 ( .A(KEYINPUT41), .ZN(n436) );
  NOR2_X1 U503 ( .A1(n706), .A2(n707), .ZN(n610) );
  AND2_X1 U504 ( .A1(n350), .A2(n356), .ZN(n410) );
  AND2_X1 U505 ( .A1(n601), .A2(n353), .ZN(n471) );
  XNOR2_X1 U506 ( .A(n571), .B(n570), .ZN(n587) );
  INV_X1 U507 ( .A(G217), .ZN(n369) );
  XNOR2_X1 U508 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U509 ( .A1(n374), .A2(n370), .ZN(n649) );
  INV_X1 U510 ( .A(G210), .ZN(n371) );
  AND2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n453), .A2(n451), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n590), .B(KEYINPUT31), .ZN(n672) );
  XNOR2_X1 U514 ( .A(n736), .B(n420), .ZN(n738) );
  XNOR2_X1 U515 ( .A(n737), .B(KEYINPUT120), .ZN(n420) );
  INV_X1 U516 ( .A(n440), .ZN(n674) );
  XOR2_X1 U517 ( .A(n615), .B(n614), .Z(n350) );
  XOR2_X1 U518 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n351) );
  AND2_X1 U519 ( .A1(n445), .A2(n544), .ZN(n352) );
  AND2_X1 U520 ( .A1(n597), .A2(n596), .ZN(n353) );
  AND2_X1 U521 ( .A1(n350), .A2(n430), .ZN(n354) );
  AND2_X1 U522 ( .A1(n686), .A2(n417), .ZN(n355) );
  AND2_X1 U523 ( .A1(n430), .A2(n408), .ZN(n356) );
  XNOR2_X1 U524 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n357) );
  XOR2_X1 U525 ( .A(KEYINPUT36), .B(KEYINPUT111), .Z(n358) );
  XOR2_X1 U526 ( .A(n529), .B(KEYINPUT104), .Z(n359) );
  INV_X1 U527 ( .A(n578), .ZN(n458) );
  XNOR2_X1 U528 ( .A(n577), .B(KEYINPUT66), .ZN(n578) );
  XNOR2_X1 U529 ( .A(n648), .B(n647), .ZN(n360) );
  XNOR2_X1 U530 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  INV_X1 U531 ( .A(n640), .ZN(n544) );
  XNOR2_X1 U532 ( .A(KEYINPUT46), .B(KEYINPUT89), .ZN(n361) );
  INV_X1 U533 ( .A(KEYINPUT45), .ZN(n485) );
  NOR2_X1 U534 ( .A1(n441), .A2(G952), .ZN(n739) );
  INV_X1 U535 ( .A(n739), .ZN(n437) );
  XOR2_X1 U536 ( .A(KEYINPUT88), .B(KEYINPUT56), .Z(n362) );
  INV_X1 U537 ( .A(G953), .ZN(n684) );
  INV_X1 U538 ( .A(n582), .ZN(n363) );
  NAND2_X1 U539 ( .A1(n366), .A2(n364), .ZN(n393) );
  NAND2_X1 U540 ( .A1(n367), .A2(n388), .ZN(n366) );
  NOR2_X1 U541 ( .A1(n643), .A2(n681), .ZN(n376) );
  NAND2_X1 U542 ( .A1(n374), .A2(n368), .ZN(n645) );
  NOR2_X1 U543 ( .A1(n681), .A2(n369), .ZN(n368) );
  NOR2_X1 U544 ( .A1(n681), .A2(n371), .ZN(n370) );
  NAND2_X1 U545 ( .A1(n374), .A2(n372), .ZN(n732) );
  NOR2_X1 U546 ( .A1(n681), .A2(n375), .ZN(n372) );
  NAND2_X1 U547 ( .A1(n374), .A2(n373), .ZN(n652) );
  NOR2_X1 U548 ( .A1(n681), .A2(n528), .ZN(n373) );
  INV_X1 U549 ( .A(n643), .ZN(n374) );
  NAND2_X1 U550 ( .A1(n376), .A2(G469), .ZN(n726) );
  NAND2_X1 U551 ( .A1(n376), .A2(G478), .ZN(n736) );
  INV_X1 U552 ( .A(n604), .ZN(n378) );
  XNOR2_X1 U553 ( .A(n489), .B(n379), .ZN(n604) );
  NAND2_X1 U554 ( .A1(n382), .A2(n461), .ZN(n460) );
  NAND2_X1 U555 ( .A1(n618), .A2(n382), .ZN(n381) );
  XNOR2_X2 U556 ( .A(n547), .B(KEYINPUT19), .ZN(n382) );
  NOR2_X1 U557 ( .A1(n676), .A2(n383), .ZN(n641) );
  XNOR2_X2 U558 ( .A(n389), .B(n485), .ZN(n383) );
  INV_X1 U559 ( .A(n383), .ZN(n384) );
  NAND2_X1 U560 ( .A1(n383), .A2(n468), .ZN(n445) );
  NAND2_X1 U561 ( .A1(n383), .A2(n678), .ZN(n679) );
  AND2_X1 U562 ( .A1(n384), .A2(n684), .ZN(n745) );
  AND2_X1 U563 ( .A1(n398), .A2(n355), .ZN(n397) );
  NAND2_X1 U564 ( .A1(n769), .A2(n765), .ZN(n464) );
  NAND2_X1 U565 ( .A1(n463), .A2(n465), .ZN(n386) );
  XNOR2_X1 U566 ( .A(n387), .B(n510), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n393), .A2(n390), .ZN(n389) );
  NAND2_X1 U568 ( .A1(n434), .A2(n433), .ZN(n392) );
  NAND2_X1 U569 ( .A1(n394), .A2(n415), .ZN(n573) );
  NAND2_X1 U570 ( .A1(n396), .A2(n628), .ZN(n395) );
  NAND2_X1 U571 ( .A1(n398), .A2(n691), .ZN(n591) );
  OR2_X1 U572 ( .A1(n650), .A2(n403), .ZN(n402) );
  NAND2_X1 U573 ( .A1(n650), .A2(G472), .ZN(n407) );
  INV_X1 U574 ( .A(n634), .ZN(n408) );
  XNOR2_X2 U575 ( .A(G113), .B(KEYINPUT3), .ZN(n413) );
  NAND2_X1 U576 ( .A1(n697), .A2(n414), .ZN(n590) );
  XNOR2_X2 U577 ( .A(n460), .B(n357), .ZN(n414) );
  INV_X1 U578 ( .A(n686), .ZN(n416) );
  INV_X1 U579 ( .A(KEYINPUT34), .ZN(n417) );
  INV_X1 U580 ( .A(KEYINPUT95), .ZN(n418) );
  INV_X1 U581 ( .A(n672), .ZN(n429) );
  XNOR2_X1 U582 ( .A(n610), .B(n436), .ZN(n700) );
  XNOR2_X1 U583 ( .A(n464), .B(n361), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n753), .B(n503), .ZN(n723) );
  XNOR2_X1 U585 ( .A(n421), .B(n362), .ZN(G51) );
  NAND2_X1 U586 ( .A1(n438), .A2(n437), .ZN(n421) );
  XNOR2_X1 U587 ( .A(n422), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U588 ( .A1(n423), .A2(n437), .ZN(n422) );
  XNOR2_X1 U589 ( .A(n645), .B(n424), .ZN(n423) );
  INV_X1 U590 ( .A(n644), .ZN(n424) );
  NAND2_X1 U591 ( .A1(n457), .A2(n578), .ZN(n456) );
  NAND2_X1 U592 ( .A1(n427), .A2(n435), .ZN(n434) );
  NAND2_X1 U593 ( .A1(n429), .A2(n428), .ZN(n427) );
  NOR2_X1 U594 ( .A1(n763), .A2(KEYINPUT87), .ZN(n483) );
  NAND2_X1 U595 ( .A1(n666), .A2(n622), .ZN(n432) );
  INV_X1 U596 ( .A(n655), .ZN(n433) );
  INV_X1 U597 ( .A(n708), .ZN(n435) );
  NAND2_X1 U598 ( .A1(n676), .A2(n468), .ZN(n467) );
  NAND2_X1 U599 ( .A1(n700), .A2(n618), .ZN(n612) );
  XNOR2_X1 U600 ( .A(n649), .B(n360), .ZN(n438) );
  NAND2_X1 U601 ( .A1(n638), .A2(n668), .ZN(n603) );
  XNOR2_X1 U602 ( .A(n602), .B(KEYINPUT39), .ZN(n638) );
  XNOR2_X1 U603 ( .A(n444), .B(n654), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n580), .A2(n578), .ZN(n455) );
  XNOR2_X2 U605 ( .A(n574), .B(n575), .ZN(n580) );
  NOR2_X1 U606 ( .A1(n580), .A2(n576), .ZN(n583) );
  NAND2_X1 U607 ( .A1(n613), .A2(n458), .ZN(n452) );
  INV_X1 U608 ( .A(n580), .ZN(n453) );
  INV_X1 U609 ( .A(KEYINPUT2), .ZN(n468) );
  NAND2_X1 U610 ( .A1(n443), .A2(n692), .ZN(n693) );
  NAND2_X1 U611 ( .A1(n443), .A2(n691), .ZN(n579) );
  NAND2_X1 U612 ( .A1(n354), .A2(n443), .ZN(n633) );
  NAND2_X1 U613 ( .A1(n583), .A2(n443), .ZN(n584) );
  NAND2_X2 U614 ( .A1(n479), .A2(n478), .ZN(n676) );
  AND2_X2 U615 ( .A1(n480), .A2(n481), .ZN(n479) );
  NAND2_X1 U616 ( .A1(n637), .A2(n484), .ZN(n480) );
  AND2_X1 U617 ( .A1(n763), .A2(KEYINPUT87), .ZN(n484) );
  NAND2_X1 U618 ( .A1(n553), .A2(G221), .ZN(n512) );
  NAND2_X1 U619 ( .A1(n506), .A2(G234), .ZN(n487) );
  XNOR2_X2 U620 ( .A(n518), .B(n517), .ZN(n687) );
  XNOR2_X2 U621 ( .A(n642), .B(KEYINPUT75), .ZN(n681) );
  XNOR2_X1 U622 ( .A(KEYINPUT94), .B(n537), .ZN(n492) );
  NAND2_X1 U623 ( .A1(G210), .A2(n546), .ZN(n493) );
  XOR2_X1 U624 ( .A(n498), .B(n497), .Z(n494) );
  AND2_X1 U625 ( .A1(n665), .A2(n631), .ZN(n495) );
  INV_X1 U626 ( .A(KEYINPUT106), .ZN(n614) );
  INV_X1 U627 ( .A(G472), .ZN(n528) );
  XNOR2_X1 U628 ( .A(n540), .B(n525), .ZN(n526) );
  XNOR2_X1 U629 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n527), .B(n526), .ZN(n650) );
  XNOR2_X1 U631 ( .A(n605), .B(KEYINPUT28), .ZN(n608) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(G475), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U634 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U635 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n611) );
  XNOR2_X1 U636 ( .A(n612), .B(n611), .ZN(n765) );
  NAND2_X1 U637 ( .A1(G227), .A2(n441), .ZN(n499) );
  XNOR2_X1 U638 ( .A(n740), .B(KEYINPUT73), .ZN(n500) );
  XOR2_X1 U639 ( .A(KEYINPUT68), .B(G101), .Z(n522) );
  INV_X1 U640 ( .A(n534), .ZN(n501) );
  NOR2_X1 U641 ( .A1(n723), .A2(G902), .ZN(n504) );
  XNOR2_X2 U642 ( .A(n504), .B(G469), .ZN(n606) );
  XNOR2_X1 U643 ( .A(n505), .B(G140), .ZN(n754) );
  XOR2_X1 U644 ( .A(G146), .B(n754), .Z(n563) );
  XOR2_X1 U645 ( .A(G137), .B(G119), .Z(n508) );
  XNOR2_X1 U646 ( .A(G128), .B(G110), .ZN(n507) );
  XNOR2_X1 U647 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U648 ( .A(n511), .B(n512), .ZN(n513) );
  XOR2_X1 U649 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n516) );
  NAND2_X1 U650 ( .A1(G234), .A2(n640), .ZN(n514) );
  NAND2_X1 U651 ( .A1(n519), .A2(G217), .ZN(n515) );
  XNOR2_X1 U652 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U653 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n520) );
  NAND2_X1 U654 ( .A1(n687), .A2(n688), .ZN(n521) );
  XOR2_X1 U655 ( .A(n522), .B(KEYINPUT5), .Z(n524) );
  NAND2_X1 U656 ( .A1(n565), .A2(G210), .ZN(n523) );
  XNOR2_X1 U657 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U658 ( .A(KEYINPUT33), .B(KEYINPUT92), .Z(n529) );
  XNOR2_X1 U659 ( .A(n531), .B(KEYINPUT14), .ZN(n597) );
  INV_X1 U660 ( .A(n597), .ZN(n716) );
  NOR2_X1 U661 ( .A1(G898), .A2(n684), .ZN(n743) );
  NAND2_X1 U662 ( .A1(n743), .A2(G902), .ZN(n532) );
  NAND2_X1 U663 ( .A1(G952), .A2(n684), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n532), .A2(n594), .ZN(n548) );
  NAND2_X1 U665 ( .A1(G224), .A2(n441), .ZN(n535) );
  XNOR2_X1 U666 ( .A(G122), .B(G104), .ZN(n564) );
  XNOR2_X1 U667 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U668 ( .A1(n626), .A2(n703), .ZN(n547) );
  XNOR2_X1 U669 ( .A(KEYINPUT101), .B(G478), .ZN(n559) );
  XOR2_X1 U670 ( .A(KEYINPUT9), .B(G122), .Z(n550) );
  XNOR2_X1 U671 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U672 ( .A(n552), .B(n551), .ZN(n557) );
  XOR2_X1 U673 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n555) );
  NAND2_X1 U674 ( .A1(G217), .A2(n553), .ZN(n554) );
  XNOR2_X1 U675 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U676 ( .A(n557), .B(n556), .ZN(n737) );
  NOR2_X1 U677 ( .A1(G902), .A2(n737), .ZN(n558) );
  XNOR2_X1 U678 ( .A(n559), .B(n558), .ZN(n586) );
  XNOR2_X1 U679 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U680 ( .A(n563), .B(n562), .Z(n569) );
  XNOR2_X1 U681 ( .A(KEYINPUT12), .B(n564), .ZN(n567) );
  NAND2_X1 U682 ( .A1(n565), .A2(G214), .ZN(n566) );
  NOR2_X1 U683 ( .A1(G902), .A2(n730), .ZN(n571) );
  NAND2_X1 U684 ( .A1(n586), .A2(n587), .ZN(n572) );
  XNOR2_X1 U685 ( .A(n572), .B(KEYINPUT105), .ZN(n628) );
  INV_X1 U686 ( .A(KEYINPUT22), .ZN(n575) );
  NOR2_X1 U687 ( .A1(n587), .A2(n586), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n577) );
  INV_X1 U689 ( .A(n687), .ZN(n585) );
  INV_X1 U690 ( .A(n598), .ZN(n691) );
  NOR2_X1 U691 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U692 ( .A1(n585), .A2(n581), .ZN(n662) );
  NAND2_X1 U693 ( .A1(n767), .A2(n662), .ZN(n582) );
  NOR2_X1 U694 ( .A1(n585), .A2(n584), .ZN(n655) );
  INV_X1 U695 ( .A(n586), .ZN(n588) );
  NOR2_X1 U696 ( .A1(n588), .A2(n587), .ZN(n671) );
  NAND2_X1 U697 ( .A1(n588), .A2(n587), .ZN(n616) );
  INV_X1 U698 ( .A(n601), .ZN(n592) );
  NOR2_X1 U699 ( .A1(n441), .A2(G900), .ZN(n593) );
  NAND2_X1 U700 ( .A1(G902), .A2(n593), .ZN(n595) );
  NAND2_X1 U701 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U702 ( .A1(n598), .A2(n703), .ZN(n599) );
  XOR2_X1 U703 ( .A(KEYINPUT30), .B(n599), .Z(n600) );
  NAND2_X1 U704 ( .A1(n625), .A2(n704), .ZN(n602) );
  NAND2_X1 U705 ( .A1(n604), .A2(n598), .ZN(n605) );
  XOR2_X1 U706 ( .A(n606), .B(KEYINPUT109), .Z(n607) );
  INV_X1 U707 ( .A(n609), .ZN(n706) );
  NAND2_X1 U708 ( .A1(n704), .A2(n703), .ZN(n707) );
  INV_X1 U709 ( .A(KEYINPUT47), .ZN(n621) );
  NOR2_X1 U710 ( .A1(KEYINPUT83), .A2(n666), .ZN(n619) );
  NOR2_X1 U711 ( .A1(n619), .A2(n708), .ZN(n620) );
  NOR2_X1 U712 ( .A1(n621), .A2(n620), .ZN(n624) );
  NOR2_X1 U713 ( .A1(KEYINPUT47), .A2(n708), .ZN(n622) );
  NOR2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n632) );
  AND2_X1 U715 ( .A1(n625), .A2(n408), .ZN(n627) );
  XNOR2_X1 U716 ( .A(KEYINPUT108), .B(n627), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n629), .A2(n628), .ZN(n665) );
  NAND2_X1 U718 ( .A1(KEYINPUT47), .A2(n381), .ZN(n630) );
  NAND2_X1 U719 ( .A1(KEYINPUT83), .A2(n630), .ZN(n631) );
  XNOR2_X1 U720 ( .A(n633), .B(KEYINPUT43), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U722 ( .A(KEYINPUT107), .B(n636), .Z(n763) );
  AND2_X1 U723 ( .A1(n638), .A2(n671), .ZN(n639) );
  XOR2_X1 U724 ( .A(KEYINPUT112), .B(n639), .Z(n770) );
  NAND2_X1 U725 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  XOR2_X1 U726 ( .A(KEYINPUT91), .B(KEYINPUT55), .Z(n648) );
  XNOR2_X1 U727 ( .A(n646), .B(KEYINPUT54), .ZN(n647) );
  INV_X1 U728 ( .A(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n650), .B(KEYINPUT62), .ZN(n651) );
  XOR2_X1 U730 ( .A(G101), .B(n655), .Z(G3) );
  NAND2_X1 U731 ( .A1(n657), .A2(n668), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n656), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n659) );
  NAND2_X1 U734 ( .A1(n657), .A2(n671), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n661) );
  XOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .Z(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(G9) );
  XNOR2_X1 U738 ( .A(G110), .B(n662), .ZN(G12) );
  XOR2_X1 U739 ( .A(G128), .B(KEYINPUT29), .Z(n664) );
  NAND2_X1 U740 ( .A1(n666), .A2(n671), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n664), .B(n663), .ZN(G30) );
  XNOR2_X1 U742 ( .A(G143), .B(n665), .ZN(G45) );
  NAND2_X1 U743 ( .A1(n666), .A2(n668), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n667), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n672), .A2(n668), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(KEYINPUT114), .ZN(n670) );
  XNOR2_X1 U747 ( .A(G113), .B(n670), .ZN(G15) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n673), .B(G116), .ZN(G18) );
  XNOR2_X1 U750 ( .A(n674), .B(G125), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n675), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U752 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n678) );
  NAND2_X1 U753 ( .A1(n678), .A2(n676), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT86), .ZN(n683) );
  XNOR2_X1 U755 ( .A(KEYINPUT85), .B(n679), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U758 ( .A1(n685), .A2(n684), .ZN(n721) );
  NAND2_X1 U759 ( .A1(n686), .A2(n700), .ZN(n719) );
  NOR2_X1 U760 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U761 ( .A(n689), .B(KEYINPUT49), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT50), .B(n693), .Z(n694) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U766 ( .A(KEYINPUT115), .B(n698), .Z(n699) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n699), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U769 ( .A(KEYINPUT116), .B(n702), .Z(n713) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n711), .A2(n416), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n717), .A2(G952), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n722), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n725) );
  XNOR2_X1 U783 ( .A(n723), .B(KEYINPUT117), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n725), .B(n724), .ZN(n727) );
  XOR2_X1 U785 ( .A(n727), .B(n726), .Z(n728) );
  NOR2_X1 U786 ( .A1(n739), .A2(n728), .ZN(G54) );
  XOR2_X1 U787 ( .A(KEYINPUT118), .B(KEYINPUT59), .Z(n729) );
  XOR2_X1 U788 ( .A(KEYINPUT60), .B(KEYINPUT119), .Z(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(G60) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(G63) );
  XNOR2_X1 U791 ( .A(n740), .B(G101), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n744) );
  NOR2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n752) );
  XNOR2_X1 U794 ( .A(n745), .B(KEYINPUT123), .ZN(n750) );
  NAND2_X1 U795 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n746), .B(KEYINPUT61), .ZN(n747) );
  XNOR2_X1 U797 ( .A(KEYINPUT122), .B(n747), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(G69) );
  XOR2_X1 U801 ( .A(n753), .B(n754), .Z(n758) );
  XNOR2_X1 U802 ( .A(G227), .B(n758), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(G953), .ZN(n757) );
  XOR2_X1 U805 ( .A(KEYINPUT125), .B(n757), .Z(n762) );
  XNOR2_X1 U806 ( .A(n676), .B(n758), .ZN(n759) );
  XNOR2_X1 U807 ( .A(n759), .B(KEYINPUT124), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(n441), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U810 ( .A(G140), .B(n763), .ZN(G42) );
  XOR2_X1 U811 ( .A(G137), .B(KEYINPUT127), .Z(n764) );
  XNOR2_X1 U812 ( .A(n765), .B(n764), .ZN(G39) );
  XOR2_X1 U813 ( .A(n766), .B(G122), .Z(G24) );
  XNOR2_X1 U814 ( .A(n767), .B(G119), .ZN(n768) );
  XNOR2_X1 U815 ( .A(n768), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U816 ( .A(G131), .B(n769), .ZN(G33) );
  XNOR2_X1 U817 ( .A(G134), .B(n770), .ZN(G36) );
endmodule

