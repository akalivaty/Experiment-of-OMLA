

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U557 ( .A1(n541), .A2(G2104), .ZN(n879) );
  XNOR2_X1 U558 ( .A(n668), .B(KEYINPUT31), .ZN(n669) );
  INV_X1 U559 ( .A(KEYINPUT96), .ZN(n668) );
  NOR2_X2 U560 ( .A1(n596), .A2(n712), .ZN(n644) );
  INV_X1 U561 ( .A(n644), .ZN(n659) );
  AND2_X1 U562 ( .A1(n700), .A2(n708), .ZN(n524) );
  NOR2_X1 U563 ( .A1(n708), .A2(n691), .ZN(n525) );
  XNOR2_X2 U564 ( .A(n554), .B(KEYINPUT65), .ZN(G160) );
  XNOR2_X1 U565 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U566 ( .A(G651), .ZN(n527) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  OR2_X1 U568 ( .A1(n527), .A2(n577), .ZN(n526) );
  XNOR2_X1 U569 ( .A(KEYINPUT67), .B(n526), .ZN(n791) );
  NAND2_X1 U570 ( .A1(G75), .A2(n791), .ZN(n536) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n787) );
  NAND2_X1 U572 ( .A1(G88), .A2(n787), .ZN(n530) );
  NOR2_X1 U573 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n528), .Z(n788) );
  NAND2_X1 U575 ( .A1(G62), .A2(n788), .ZN(n529) );
  NAND2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n534) );
  NOR2_X1 U577 ( .A1(G651), .A2(n577), .ZN(n531) );
  XNOR2_X1 U578 ( .A(KEYINPUT64), .B(n531), .ZN(n792) );
  NAND2_X1 U579 ( .A1(n792), .A2(G50), .ZN(n532) );
  XOR2_X1 U580 ( .A(KEYINPUT80), .B(n532), .Z(n533) );
  NOR2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U583 ( .A(n537), .B(KEYINPUT81), .Z(G303) );
  INV_X1 U584 ( .A(G303), .ZN(G166) );
  INV_X1 U585 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U586 ( .A1(G102), .A2(n879), .ZN(n540) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n538), .Z(n719) );
  NAND2_X1 U589 ( .A1(G138), .A2(n719), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n546) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U592 ( .A1(G114), .A2(n883), .ZN(n544) );
  NOR2_X1 U593 ( .A1(n541), .A2(G2104), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT66), .ZN(n715) );
  NAND2_X1 U595 ( .A1(G126), .A2(n715), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U597 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U598 ( .A1(n715), .A2(G125), .ZN(n553) );
  NAND2_X1 U599 ( .A1(G137), .A2(n719), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G113), .A2(n883), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G101), .A2(n879), .ZN(n549) );
  XNOR2_X1 U603 ( .A(KEYINPUT23), .B(n549), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G90), .A2(n787), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G77), .A2(n791), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U609 ( .A(KEYINPUT9), .B(n557), .ZN(n561) );
  NAND2_X1 U610 ( .A1(n792), .A2(G52), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n788), .A2(G64), .ZN(n558) );
  AND2_X1 U612 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n561), .A2(n560), .ZN(G301) );
  INV_X1 U614 ( .A(G301), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n787), .A2(G89), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT4), .B(n562), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n791), .A2(G76), .ZN(n563) );
  XOR2_X1 U618 ( .A(KEYINPUT75), .B(n563), .Z(n564) );
  NAND2_X1 U619 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U620 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U621 ( .A1(n788), .A2(G63), .ZN(n568) );
  NAND2_X1 U622 ( .A1(G51), .A2(n792), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U626 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G651), .A2(G74), .ZN(n573) );
  XOR2_X1 U629 ( .A(KEYINPUT77), .B(n573), .Z(n575) );
  NAND2_X1 U630 ( .A1(G49), .A2(n792), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U632 ( .A(KEYINPUT78), .B(n576), .Z(n579) );
  NAND2_X1 U633 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U635 ( .A1(n788), .A2(n580), .ZN(n581) );
  XNOR2_X1 U636 ( .A(KEYINPUT79), .B(n581), .ZN(G288) );
  NAND2_X1 U637 ( .A1(G86), .A2(n787), .ZN(n583) );
  NAND2_X1 U638 ( .A1(G48), .A2(n792), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n791), .A2(G73), .ZN(n584) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U643 ( .A1(n788), .A2(G61), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G85), .A2(n787), .ZN(n590) );
  NAND2_X1 U646 ( .A1(G47), .A2(n792), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U648 ( .A1(G72), .A2(n791), .ZN(n591) );
  XOR2_X1 U649 ( .A(KEYINPUT68), .B(n591), .Z(n592) );
  NOR2_X1 U650 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U651 ( .A1(n788), .A2(G60), .ZN(n594) );
  NAND2_X1 U652 ( .A1(n595), .A2(n594), .ZN(G290) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n713) );
  INV_X1 U654 ( .A(n713), .ZN(n596) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n712) );
  NOR2_X1 U656 ( .A1(G2090), .A2(n659), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G8), .A2(n659), .ZN(n708) );
  NOR2_X1 U658 ( .A1(G1971), .A2(n708), .ZN(n597) );
  NOR2_X1 U659 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U660 ( .A(KEYINPUT98), .B(n599), .Z(n600) );
  NOR2_X1 U661 ( .A1(G166), .A2(n600), .ZN(n601) );
  XNOR2_X1 U662 ( .A(KEYINPUT99), .B(n601), .ZN(n675) );
  INV_X1 U663 ( .A(G1961), .ZN(n832) );
  NAND2_X1 U664 ( .A1(n659), .A2(n832), .ZN(n604) );
  XOR2_X1 U665 ( .A(G2078), .B(KEYINPUT93), .Z(n602) );
  XNOR2_X1 U666 ( .A(KEYINPUT25), .B(n602), .ZN(n1014) );
  NAND2_X1 U667 ( .A1(n644), .A2(n1014), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n665) );
  NAND2_X1 U669 ( .A1(n665), .A2(G171), .ZN(n658) );
  NAND2_X1 U670 ( .A1(n644), .A2(G2072), .ZN(n605) );
  XNOR2_X1 U671 ( .A(n605), .B(KEYINPUT27), .ZN(n607) );
  AND2_X1 U672 ( .A1(G1956), .A2(n659), .ZN(n606) );
  NOR2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n616) );
  NAND2_X1 U674 ( .A1(n788), .A2(G65), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G53), .A2(n792), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G91), .A2(n787), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G78), .A2(n791), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n983) );
  NOR2_X1 U681 ( .A1(n616), .A2(n983), .ZN(n615) );
  XOR2_X1 U682 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n614) );
  XNOR2_X1 U683 ( .A(n615), .B(n614), .ZN(n655) );
  NAND2_X1 U684 ( .A1(n616), .A2(n983), .ZN(n653) );
  XOR2_X1 U685 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n618) );
  NAND2_X1 U686 ( .A1(G56), .A2(n788), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(n625) );
  NAND2_X1 U688 ( .A1(G81), .A2(n787), .ZN(n619) );
  XOR2_X1 U689 ( .A(KEYINPUT12), .B(n619), .Z(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT73), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G68), .A2(n791), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U693 ( .A(KEYINPUT13), .B(n623), .Z(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G43), .A2(n792), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n989) );
  INV_X1 U697 ( .A(G1341), .ZN(n990) );
  NOR2_X1 U698 ( .A1(n644), .A2(n990), .ZN(n628) );
  NAND2_X1 U699 ( .A1(KEYINPUT26), .A2(n628), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n630), .A2(KEYINPUT95), .ZN(n635) );
  INV_X1 U701 ( .A(KEYINPUT95), .ZN(n633) );
  NAND2_X1 U702 ( .A1(G1996), .A2(n644), .ZN(n629) );
  XNOR2_X1 U703 ( .A(KEYINPUT26), .B(n629), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n989), .A2(n636), .ZN(n648) );
  NAND2_X1 U708 ( .A1(n791), .A2(G79), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G54), .A2(n792), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G92), .A2(n787), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G66), .A2(n788), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U715 ( .A(n643), .B(KEYINPUT15), .Z(n978) );
  INV_X1 U716 ( .A(n978), .ZN(n768) );
  NAND2_X1 U717 ( .A1(G1348), .A2(n659), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G2067), .A2(n644), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n649) );
  NOR2_X1 U720 ( .A1(n768), .A2(n649), .ZN(n647) );
  OR2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n768), .A2(n649), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U726 ( .A(KEYINPUT29), .B(n656), .Z(n657) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n672) );
  NOR2_X1 U728 ( .A1(n659), .A2(G2084), .ZN(n660) );
  XOR2_X1 U729 ( .A(n660), .B(KEYINPUT91), .Z(n678) );
  INV_X1 U730 ( .A(G8), .ZN(n661) );
  OR2_X1 U731 ( .A1(n678), .A2(n661), .ZN(n662) );
  NOR2_X1 U732 ( .A1(G1966), .A2(n708), .ZN(n682) );
  NOR2_X1 U733 ( .A1(n662), .A2(n682), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT30), .B(n663), .Z(n664) );
  NOR2_X1 U735 ( .A1(G168), .A2(n664), .ZN(n667) );
  NOR2_X1 U736 ( .A1(G171), .A2(n665), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n680) );
  NAND2_X1 U739 ( .A1(n680), .A2(G286), .ZN(n673) );
  XOR2_X1 U740 ( .A(n673), .B(KEYINPUT97), .Z(n674) );
  NAND2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n676), .A2(G8), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n677), .B(KEYINPUT32), .ZN(n686) );
  NAND2_X1 U744 ( .A1(G8), .A2(n678), .ZN(n679) );
  XNOR2_X1 U745 ( .A(KEYINPUT92), .B(n679), .ZN(n684) );
  INV_X1 U746 ( .A(n680), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n698) );
  NOR2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NOR2_X1 U751 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n690), .A2(n687), .ZN(n998) );
  NAND2_X1 U753 ( .A1(n698), .A2(n998), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT100), .ZN(n695) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U756 ( .A(n987), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n708), .A2(n689), .ZN(n693) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n995) );
  INV_X1 U759 ( .A(n995), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n690), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U761 ( .A1(n692), .A2(n525), .ZN(n696) );
  AND2_X1 U762 ( .A1(n693), .A2(n696), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n703) );
  AND2_X1 U764 ( .A1(n696), .A2(KEYINPUT33), .ZN(n701) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U766 ( .A1(G8), .A2(n697), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U768 ( .A1(n701), .A2(n524), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n704), .B(KEYINPUT101), .ZN(n711) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT89), .B(n705), .ZN(n706) );
  XNOR2_X1 U773 ( .A(KEYINPUT24), .B(n706), .ZN(n707) );
  NOR2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U775 ( .A(KEYINPUT90), .B(n709), .Z(n710) );
  NAND2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n749) );
  XNOR2_X1 U777 ( .A(G1986), .B(G290), .ZN(n980) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U779 ( .A(KEYINPUT83), .B(n714), .ZN(n745) );
  INV_X1 U780 ( .A(n745), .ZN(n760) );
  NAND2_X1 U781 ( .A1(n980), .A2(n760), .ZN(n747) );
  NAND2_X1 U782 ( .A1(G116), .A2(n883), .ZN(n717) );
  BUF_X1 U783 ( .A(n715), .Z(n884) );
  NAND2_X1 U784 ( .A1(G128), .A2(n884), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n718), .B(KEYINPUT35), .ZN(n724) );
  NAND2_X1 U787 ( .A1(G104), .A2(n879), .ZN(n721) );
  BUF_X1 U788 ( .A(n719), .Z(n880) );
  NAND2_X1 U789 ( .A1(G140), .A2(n880), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U791 ( .A(KEYINPUT34), .B(n722), .Z(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U793 ( .A(n725), .B(KEYINPUT36), .Z(n893) );
  XNOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  OR2_X1 U795 ( .A1(n893), .A2(n758), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n726), .B(KEYINPUT84), .ZN(n930) );
  NOR2_X1 U797 ( .A1(n745), .A2(n930), .ZN(n727) );
  XOR2_X1 U798 ( .A(n727), .B(KEYINPUT85), .Z(n755) );
  XOR2_X1 U799 ( .A(KEYINPUT87), .B(G1991), .Z(n1015) );
  NAND2_X1 U800 ( .A1(G131), .A2(n880), .ZN(n729) );
  NAND2_X1 U801 ( .A1(G119), .A2(n884), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G95), .A2(n879), .ZN(n731) );
  NAND2_X1 U804 ( .A1(G107), .A2(n883), .ZN(n730) );
  NAND2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U807 ( .A(n734), .B(KEYINPUT86), .Z(n860) );
  AND2_X1 U808 ( .A1(n1015), .A2(n860), .ZN(n744) );
  XOR2_X1 U809 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n736) );
  NAND2_X1 U810 ( .A1(G105), .A2(n879), .ZN(n735) );
  XNOR2_X1 U811 ( .A(n736), .B(n735), .ZN(n740) );
  NAND2_X1 U812 ( .A1(G117), .A2(n883), .ZN(n738) );
  NAND2_X1 U813 ( .A1(G129), .A2(n884), .ZN(n737) );
  NAND2_X1 U814 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n880), .A2(G141), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n742), .A2(n741), .ZN(n863) );
  AND2_X1 U818 ( .A1(n863), .A2(G1996), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n941) );
  NOR2_X1 U820 ( .A1(n941), .A2(n745), .ZN(n752) );
  NOR2_X1 U821 ( .A1(n755), .A2(n752), .ZN(n746) );
  AND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n763) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n863), .ZN(n933) );
  NOR2_X1 U825 ( .A1(n1015), .A2(n860), .ZN(n939) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U827 ( .A1(n939), .A2(n750), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U829 ( .A1(n933), .A2(n753), .ZN(n754) );
  XNOR2_X1 U830 ( .A(n754), .B(KEYINPUT39), .ZN(n757) );
  INV_X1 U831 ( .A(n755), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n758), .A2(n893), .ZN(n942) );
  NAND2_X1 U834 ( .A1(n759), .A2(n942), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G82), .ZN(G220) );
  XOR2_X1 U841 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n766) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XOR2_X1 U843 ( .A(n766), .B(n765), .Z(n821) );
  NAND2_X1 U844 ( .A1(n821), .A2(G567), .ZN(n767) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  INV_X1 U846 ( .A(G860), .ZN(n920) );
  OR2_X1 U847 ( .A1(n989), .A2(n920), .ZN(G153) );
  INV_X1 U848 ( .A(G868), .ZN(n805) );
  NAND2_X1 U849 ( .A1(n768), .A2(n805), .ZN(n769) );
  XNOR2_X1 U850 ( .A(n769), .B(KEYINPUT74), .ZN(n771) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n770) );
  NAND2_X1 U852 ( .A1(n771), .A2(n770), .ZN(G284) );
  XNOR2_X1 U853 ( .A(n983), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U854 ( .A1(G286), .A2(G868), .ZN(n773) );
  NAND2_X1 U855 ( .A1(G299), .A2(n805), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n920), .A2(G559), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n774), .A2(n978), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n775), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n989), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G868), .A2(n978), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G99), .A2(n879), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G111), .A2(n883), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n884), .A2(G123), .ZN(n781) );
  XNOR2_X1 U868 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n880), .A2(G135), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n938) );
  XNOR2_X1 U872 ( .A(n938), .B(G2096), .ZN(n786) );
  INV_X1 U873 ( .A(G2100), .ZN(n845) );
  NAND2_X1 U874 ( .A1(n786), .A2(n845), .ZN(G156) );
  NAND2_X1 U875 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U878 ( .A1(n791), .A2(G80), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U882 ( .A(KEYINPUT76), .B(n797), .Z(n921) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(n921), .ZN(n799) );
  XOR2_X1 U884 ( .A(G305), .B(G303), .Z(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n802) );
  XNOR2_X1 U886 ( .A(G290), .B(G288), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n800), .B(G299), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n802), .B(n801), .ZN(n896) );
  NAND2_X1 U889 ( .A1(G559), .A2(n978), .ZN(n803) );
  XOR2_X1 U890 ( .A(n989), .B(n803), .Z(n919) );
  XOR2_X1 U891 ( .A(n896), .B(n919), .Z(n804) );
  NOR2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n807) );
  NOR2_X1 U893 ( .A1(n921), .A2(G868), .ZN(n806) );
  NOR2_X1 U894 ( .A1(n807), .A2(n806), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2084), .A2(G2078), .ZN(n808) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XOR2_X1 U900 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U901 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U902 ( .A1(G108), .A2(G120), .ZN(n812) );
  NOR2_X1 U903 ( .A1(G237), .A2(n812), .ZN(n813) );
  NAND2_X1 U904 ( .A1(G69), .A2(n813), .ZN(n923) );
  NAND2_X1 U905 ( .A1(n923), .A2(G567), .ZN(n818) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U908 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U909 ( .A1(G96), .A2(n816), .ZN(n924) );
  NAND2_X1 U910 ( .A1(n924), .A2(G2106), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n826) );
  NAND2_X1 U912 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n826), .A2(n819), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n825), .A2(G36), .ZN(n820) );
  XNOR2_X1 U915 ( .A(KEYINPUT82), .B(n820), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n821), .ZN(G217) );
  INV_X1 U917 ( .A(n821), .ZN(G223) );
  NAND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n822) );
  XOR2_X1 U919 ( .A(KEYINPUT104), .B(n822), .Z(n823) );
  NAND2_X1 U920 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U923 ( .A(n826), .ZN(G319) );
  XOR2_X1 U924 ( .A(KEYINPUT108), .B(G1956), .Z(n828) );
  XNOR2_X1 U925 ( .A(G1996), .B(G1991), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U927 ( .A(n829), .B(KEYINPUT107), .Z(n831) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1971), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n836) );
  XNOR2_X1 U930 ( .A(G1976), .B(n832), .ZN(n834) );
  XNOR2_X1 U931 ( .A(G1981), .B(G1966), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U934 ( .A(G2474), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2678), .Z(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2072), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n847) );
  XOR2_X1 U943 ( .A(G2096), .B(n845), .Z(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U945 ( .A(G2084), .B(G2078), .Z(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(G227) );
  NAND2_X1 U947 ( .A1(G136), .A2(n880), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT110), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G112), .A2(n883), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT111), .B(n851), .Z(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U952 ( .A1(n884), .A2(G124), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n854), .Z(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT109), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G100), .A2(n879), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U958 ( .A(n938), .B(G162), .Z(n862) );
  XNOR2_X1 U959 ( .A(G164), .B(n860), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n878) );
  XOR2_X1 U961 ( .A(n863), .B(KEYINPUT48), .Z(n876) );
  XNOR2_X1 U962 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G106), .A2(n879), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G142), .A2(n880), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT45), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G118), .A2(n883), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G130), .A2(n884), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(n878), .B(n877), .Z(n892) );
  NAND2_X1 U976 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U979 ( .A1(G115), .A2(n883), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G127), .A2(n884), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(KEYINPUT115), .B(n887), .ZN(n888) );
  XNOR2_X1 U983 ( .A(KEYINPUT47), .B(n888), .ZN(n889) );
  NOR2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n926) );
  XNOR2_X1 U985 ( .A(G160), .B(n926), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U987 ( .A(n894), .B(n893), .Z(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n896), .B(KEYINPUT116), .ZN(n898) );
  XOR2_X1 U990 ( .A(n978), .B(G286), .Z(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U992 ( .A(n989), .B(G301), .Z(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U994 ( .A1(G37), .A2(n901), .ZN(n902) );
  XOR2_X1 U995 ( .A(KEYINPUT117), .B(n902), .Z(G397) );
  XNOR2_X1 U996 ( .A(G2451), .B(G2427), .ZN(n912) );
  XOR2_X1 U997 ( .A(G2430), .B(G2443), .Z(n904) );
  XNOR2_X1 U998 ( .A(KEYINPUT103), .B(G2438), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n906) );
  XOR2_X1 U1001 ( .A(n990), .B(G1348), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1004 ( .A(G2446), .B(KEYINPUT102), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n913), .A2(G14), .ZN(n925) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n925), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  XOR2_X1 U1014 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(G145) );
  INV_X1 U1018 ( .A(G120), .ZN(G236) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(G325) );
  INV_X1 U1023 ( .A(G325), .ZN(G261) );
  INV_X1 U1024 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1025 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT50), .B(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G162), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT119), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT51), .B(n935), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n947) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G2084), .B(G160), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n948), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n949), .B(KEYINPUT120), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(KEYINPUT55), .A2(n950), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(n951), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G29), .ZN(n1008) );
  XOR2_X1 U1046 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n959) );
  XNOR2_X1 U1047 ( .A(G1986), .B(G24), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G1971), .B(G22), .Z(n955) );
  XNOR2_X1 U1051 ( .A(KEYINPUT126), .B(n955), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n959), .B(n958), .ZN(n973) );
  XOR2_X1 U1054 ( .A(G5), .B(G1961), .Z(n971) );
  XOR2_X1 U1055 ( .A(G19), .B(G1341), .Z(n963) );
  XNOR2_X1 U1056 ( .A(G1981), .B(G6), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G1956), .B(G20), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT59), .B(G1348), .Z(n964) );
  XNOR2_X1 U1061 ( .A(G4), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1063 ( .A(KEYINPUT60), .B(n967), .Z(n969) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT61), .B(n974), .ZN(n975) );
  INV_X1 U1069 ( .A(G16), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n977), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(G11), .ZN(n1006) );
  XNOR2_X1 U1072 ( .A(n977), .B(KEYINPUT56), .ZN(n1003) );
  XOR2_X1 U1073 ( .A(G1348), .B(n978), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(G1971), .A2(G303), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n986) );
  XOR2_X1 U1077 ( .A(G1956), .B(n983), .Z(n984) );
  XNOR2_X1 U1078 ( .A(KEYINPUT124), .B(n984), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n994) );
  XOR2_X1 U1080 ( .A(G301), .B(G1961), .Z(n988) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n992) );
  XOR2_X1 U1082 ( .A(n990), .B(n989), .Z(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT57), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT125), .B(n1004), .Z(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1031) );
  XOR2_X1 U1094 ( .A(G2072), .B(G33), .Z(n1009) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(G28), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(G2067), .B(G26), .Z(n1011) );
  XOR2_X1 U1097 ( .A(G1996), .B(G32), .Z(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1100 ( .A(n1014), .B(G27), .Z(n1017) );
  XNOR2_X1 U1101 ( .A(n1015), .B(G25), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(n1020), .B(KEYINPUT53), .ZN(n1023) );
  XOR2_X1 U1105 ( .A(G2084), .B(G34), .Z(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(KEYINPUT122), .B(G2090), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(G35), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT55), .B(n1027), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT123), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1113 ( .A1(G29), .A2(n1029), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(n1032), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

