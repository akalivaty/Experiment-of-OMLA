//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(G134), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G122), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G107), .B(new_n194), .C1(new_n196), .C2(KEYINPUT14), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT89), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT13), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n188), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n187), .A3(new_n206), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n202), .A2(new_n207), .B1(new_n208), .B2(new_n191), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(new_n188), .A3(KEYINPUT89), .A4(new_n206), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n199), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n195), .A2(new_n198), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n212), .A2(new_n213), .B1(G134), .B2(new_n191), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT90), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n202), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n191), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n210), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n191), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(new_n213), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n199), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT90), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n200), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT9), .B(G234), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n226), .A2(new_n227), .A3(G953), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT91), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n200), .B(new_n228), .C1(new_n216), .C2(new_n224), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  INV_X1    g049(.A(new_n200), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n215), .B1(new_n211), .B2(new_n214), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(KEYINPUT90), .A3(new_n223), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT91), .A3(new_n228), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G478), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT15), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G475), .ZN(new_n246));
  NOR2_X1   g060(.A1(G237), .A2(G953), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n247), .A2(G143), .A3(G214), .ZN(new_n248));
  AOI21_X1  g062(.A(G143), .B1(new_n247), .B2(G214), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n187), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n247), .A2(G143), .A3(G214), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n251), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G140), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  INV_X1    g075(.A(G125), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G140), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT16), .ZN(new_n264));
  OR3_X1    g078(.A1(new_n262), .A2(KEYINPUT16), .A3(G140), .ZN(new_n265));
  AOI21_X1  g079(.A(G146), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(G146), .ZN(new_n268));
  OAI211_X1 g082(.A(KEYINPUT17), .B(G131), .C1(new_n248), .C2(new_n249), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n259), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT82), .A2(KEYINPUT18), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(G131), .B(new_n272), .C1(new_n248), .C2(new_n249), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n255), .B(new_n257), .C1(new_n256), .C2(new_n271), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n263), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  INV_X1    g090(.A(G146), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n263), .A3(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n276), .A2(KEYINPUT83), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT83), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n273), .B(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(G113), .B(G122), .Z(new_n282));
  XOR2_X1   g096(.A(KEYINPUT84), .B(G104), .Z(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G113), .B(G122), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT84), .B(G104), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT85), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(new_n290), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n270), .A2(new_n281), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n270), .A2(new_n281), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n287), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n270), .B2(new_n281), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n246), .B1(new_n298), .B2(new_n235), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n301));
  NOR2_X1   g115(.A1(G475), .A2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n270), .A2(new_n281), .A3(new_n292), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n250), .A2(new_n258), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT19), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT19), .B1(new_n261), .B2(new_n263), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n277), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n268), .A2(KEYINPUT72), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n264), .A2(new_n265), .A3(new_n309), .A4(G146), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n307), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n288), .B1(new_n281), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n281), .A2(new_n311), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n293), .B1(new_n315), .B2(new_n288), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n301), .A4(new_n302), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n302), .B1(new_n303), .B2(new_n312), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n314), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n253), .A2(G952), .ZN(new_n324));
  NAND2_X1  g138(.A1(G234), .A2(G237), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT93), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT21), .B(G898), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(G902), .A3(G953), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n300), .A2(new_n323), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n241), .A2(new_n243), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n245), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G214), .B1(G237), .B2(G902), .ZN(new_n337));
  INV_X1    g151(.A(G224), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G953), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n277), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n187), .A2(G146), .ZN(new_n341));
  AOI21_X1  g155(.A(G128), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n187), .A2(KEYINPUT1), .A3(G146), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n340), .A3(new_n341), .ZN(new_n347));
  AOI21_X1  g161(.A(G125), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G143), .B(G146), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(KEYINPUT0), .A2(G128), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT0), .A2(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n340), .A2(new_n341), .A3(new_n352), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n262), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n339), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n347), .B(new_n343), .C1(G128), .C2(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n262), .ZN(new_n360));
  INV_X1    g174(.A(new_n339), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n340), .A2(new_n341), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  OAI21_X1  g176(.A(G125), .B1(new_n362), .B2(new_n355), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT7), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n358), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n360), .A2(new_n363), .A3(new_n365), .A4(new_n361), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G122), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT8), .Z(new_n371));
  INV_X1    g185(.A(G113), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT2), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G113), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G116), .B(G119), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n193), .A2(G119), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT5), .ZN(new_n382));
  OAI21_X1  g196(.A(G113), .B1(new_n380), .B2(KEYINPUT5), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n198), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n387), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n386), .A2(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n198), .A2(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n384), .A2(new_n385), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n385), .B1(new_n384), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n384), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n371), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n369), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT74), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT74), .A4(new_n391), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(G101), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n380), .A2(new_n381), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT2), .B(G113), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n378), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n418), .A3(G101), .A4(new_n410), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n404), .A3(new_n370), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n406), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n404), .ZN(new_n423));
  INV_X1    g237(.A(new_n370), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n421), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n358), .A2(new_n364), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n428), .A3(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n422), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n422), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n337), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n422), .A2(new_n430), .ZN(new_n437));
  INV_X1    g251(.A(new_n431), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n422), .A2(new_n430), .A3(new_n431), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT80), .A3(new_n337), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT75), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n342), .B2(new_n344), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT75), .B(new_n343), .C1(new_n349), .C2(G128), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n347), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n396), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g263(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n354), .A2(new_n356), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n413), .A2(new_n453), .A3(new_n419), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n201), .A2(G137), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT64), .B1(new_n456), .B2(G134), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT64), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(new_n458), .C1(new_n201), .C2(G137), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(new_n201), .B2(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n465), .A2(new_n256), .A3(new_n461), .A4(new_n455), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n401), .A2(KEYINPUT10), .A3(new_n359), .A4(new_n403), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n452), .A2(new_n454), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT12), .B1(new_n467), .B2(KEYINPUT78), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n401), .A2(new_n403), .ZN(new_n473));
  INV_X1    g287(.A(new_n359), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n448), .B2(new_n447), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n475), .B2(new_n468), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n253), .A2(G227), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n343), .B1(new_n349), .B2(G128), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(new_n444), .B1(new_n349), .B2(new_n346), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n396), .B1(new_n482), .B2(new_n446), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n359), .B1(new_n401), .B2(new_n403), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n471), .B(new_n467), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AND4_X1   g299(.A1(new_n470), .A2(new_n476), .A3(new_n480), .A4(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n469), .B1(new_n483), .B2(new_n450), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n413), .A2(new_n453), .A3(new_n419), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n480), .B1(new_n489), .B2(new_n470), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n443), .B(new_n235), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n443), .A2(new_n235), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n476), .A2(new_n470), .A3(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n479), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n470), .A3(new_n480), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(G469), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G221), .B1(new_n226), .B2(G902), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n336), .A2(new_n436), .A3(new_n442), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT70), .B1(new_n189), .B2(G119), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n379), .A3(G128), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n189), .A2(G119), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n379), .A2(G128), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n379), .A2(G128), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(KEYINPUT23), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT71), .B(G110), .Z(new_n513));
  OAI22_X1  g327(.A1(new_n507), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n308), .A3(new_n310), .A4(new_n278), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n508), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(G110), .ZN(new_n517));
  INV_X1    g331(.A(new_n268), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(new_n266), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(new_n519), .A3(new_n523), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n235), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(KEYINPUT25), .A3(new_n235), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n227), .B1(G234), .B2(new_n235), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT73), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n534));
  INV_X1    g348(.A(new_n532), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n534), .B(new_n535), .C1(new_n529), .C2(new_n530), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n515), .A2(new_n519), .A3(new_n523), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n523), .B1(new_n515), .B2(new_n519), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n532), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n416), .A2(new_n378), .A3(KEYINPUT65), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT65), .B1(new_n416), .B2(new_n378), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n463), .A2(new_n466), .B1(new_n354), .B2(new_n356), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n201), .A2(G137), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n456), .A2(G134), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n359), .A2(new_n466), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n547), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n466), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n464), .B2(KEYINPUT11), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n256), .B1(new_n555), .B2(new_n461), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n453), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT65), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n376), .A2(new_n377), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n414), .A2(new_n415), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n416), .A2(new_n378), .A3(KEYINPUT65), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n359), .A2(new_n466), .A3(new_n551), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n557), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n553), .A2(new_n565), .A3(KEYINPUT68), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT68), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n547), .B(new_n567), .C1(new_n548), .C2(new_n552), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(KEYINPUT28), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n247), .A2(G210), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT27), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT26), .B(G101), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n569), .A2(new_n571), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n581), .A2(new_n582), .A3(new_n235), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n581), .B2(new_n235), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT30), .B1(new_n548), .B2(new_n552), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT30), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n557), .A2(new_n586), .A3(new_n564), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n585), .A2(new_n587), .B1(new_n416), .B2(new_n378), .ZN(new_n588));
  INV_X1    g402(.A(new_n565), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n557), .A2(new_n563), .A3(KEYINPUT28), .A4(new_n564), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n417), .B1(new_n548), .B2(new_n552), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n576), .A2(KEYINPUT66), .A3(new_n577), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT66), .B1(new_n576), .B2(new_n577), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n571), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n590), .A2(new_n597), .A3(new_n579), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n583), .A2(new_n584), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT32), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n593), .B2(new_n571), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n548), .A2(new_n552), .A3(KEYINPUT30), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n586), .B1(new_n557), .B2(new_n564), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n417), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n578), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n565), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT31), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n585), .A2(new_n587), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n589), .B1(new_n611), .B2(new_n417), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT31), .A3(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n603), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT67), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n602), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n603), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT31), .B1(new_n612), .B2(new_n607), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n588), .A2(new_n609), .A3(new_n589), .A4(new_n578), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(KEYINPUT32), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n544), .B1(new_n601), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n502), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n390), .ZN(G3));
  OAI21_X1  g441(.A(G472), .B1(new_n614), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n622), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n630), .A2(new_n544), .A3(new_n501), .A4(KEYINPUT94), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n537), .A3(new_n629), .A4(new_n542), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n500), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT95), .B1(new_n239), .B2(new_n228), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n239), .A2(new_n228), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT33), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n232), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n230), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n636), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n641), .B2(new_n230), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(KEYINPUT96), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n233), .A2(new_n644), .A3(new_n240), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n242), .A2(G902), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n643), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n233), .A2(new_n235), .A3(new_n240), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n242), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n313), .A2(KEYINPUT86), .B1(new_n319), .B2(new_n321), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n299), .B1(new_n318), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n434), .A3(new_n332), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n635), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n322), .B2(KEYINPUT97), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n664), .B(KEYINPUT98), .C1(new_n319), .C2(new_n321), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n319), .A2(new_n321), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n666), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n320), .B1(new_n316), .B2(new_n302), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT98), .B1(new_n669), .B2(new_n664), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n322), .A2(KEYINPUT97), .A3(new_n662), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n300), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n243), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n241), .B(new_n674), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n673), .A2(new_n675), .A3(new_n434), .A4(new_n332), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n635), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n524), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n520), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n541), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n533), .A2(new_n536), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n630), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n502), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NOR3_X1   g503(.A1(new_n614), .A2(new_n602), .A3(new_n616), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT32), .B1(new_n621), .B2(new_n622), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n584), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n581), .A2(new_n582), .A3(new_n235), .ZN(new_n694));
  INV_X1    g508(.A(new_n598), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n684), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n670), .A2(new_n668), .A3(new_n671), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n299), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n241), .A2(new_n243), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n244), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n327), .B1(G900), .B2(new_n330), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n500), .A2(new_n434), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n698), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XNOR2_X1  g522(.A(new_n704), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n501), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT40), .Z(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n441), .B(new_n712), .Z(new_n713));
  INV_X1    g527(.A(new_n337), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n703), .A2(new_n656), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n713), .A2(new_n714), .A3(new_n685), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n566), .A2(new_n568), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n608), .B1(new_n596), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n235), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G472), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n617), .A2(new_n623), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n617), .A2(new_n623), .A3(new_n723), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n711), .A2(new_n716), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  INV_X1    g541(.A(new_n704), .ZN(new_n728));
  AOI211_X1 g542(.A(new_n655), .B(new_n728), .C1(new_n650), .C2(new_n652), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n698), .A2(new_n706), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  AOI21_X1  g545(.A(new_n543), .B1(new_n692), .B2(new_n697), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n235), .B1(new_n486), .B2(new_n490), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n734), .A2(new_n499), .A3(new_n491), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n658), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n676), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  INV_X1    g556(.A(KEYINPUT102), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n714), .B1(new_n439), .B2(new_n440), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n735), .A2(new_n744), .A3(KEYINPUT101), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT101), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n734), .A2(new_n499), .A3(new_n491), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n434), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n692), .A2(new_n697), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n336), .A3(new_n685), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n745), .A2(new_n748), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT102), .A3(new_n698), .A4(new_n336), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n621), .A2(new_n235), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n569), .A2(new_n571), .ZN(new_n758));
  OAI22_X1  g572(.A1(new_n758), .A2(new_n596), .B1(new_n619), .B2(new_n620), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n757), .A2(G472), .B1(new_n622), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n544), .A2(new_n333), .A3(new_n760), .A4(new_n735), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n703), .A2(new_n744), .A3(new_n656), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(G122), .Z(G24));
  NAND2_X1  g578(.A1(new_n759), .A2(new_n622), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n628), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n684), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n729), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  OAI22_X1  g584(.A1(new_n599), .A2(new_n600), .B1(new_n691), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT105), .B1(new_n617), .B2(new_n623), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n544), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT106), .B(new_n544), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n439), .A2(new_n337), .A3(new_n440), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT103), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n494), .A2(new_n779), .A3(new_n479), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n496), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n494), .B2(new_n479), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n443), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n491), .A2(new_n493), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n499), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n778), .B1(new_n785), .B2(KEYINPUT104), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n499), .C1(new_n783), .C2(new_n784), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n729), .A3(KEYINPUT42), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n732), .A2(new_n786), .A3(new_n729), .A4(new_n788), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NAND4_X1  g610(.A1(new_n732), .A2(new_n705), .A3(new_n786), .A4(new_n788), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NOR2_X1   g612(.A1(new_n781), .A2(new_n782), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n495), .B2(new_n496), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n443), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n492), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n491), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n499), .B(new_n709), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT107), .Z(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n653), .A2(new_n655), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n630), .A2(new_n684), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n778), .B1(new_n813), .B2(KEYINPUT44), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n808), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT108), .B(G137), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G39));
  OAI21_X1  g632(.A(new_n499), .B1(new_n804), .B2(new_n805), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n750), .A2(new_n544), .A3(new_n778), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n729), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n702), .A2(new_n244), .A3(new_n704), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT111), .B1(new_n673), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n500), .A2(new_n778), .A3(new_n684), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n701), .A2(new_n675), .A3(new_n831), .A4(new_n704), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .A4(new_n750), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n786), .A2(new_n729), .A3(new_n767), .A4(new_n788), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n797), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n791), .B2(new_n794), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n502), .A2(new_n625), .B1(new_n761), .B2(new_n762), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n687), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n737), .B1(new_n658), .B2(new_n676), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT109), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n657), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n653), .A2(KEYINPUT109), .A3(new_n656), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n703), .A2(new_n844), .A3(new_n655), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT110), .B1(new_n675), .B2(new_n656), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n436), .A2(new_n442), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n635), .A2(new_n847), .A3(new_n848), .A4(new_n333), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n836), .A2(new_n840), .A3(new_n755), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n851));
  INV_X1    g665(.A(new_n762), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n725), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n704), .B(KEYINPUT112), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n537), .A2(new_n854), .A3(new_n682), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT25), .B1(new_n540), .B2(new_n235), .ZN(new_n857));
  INV_X1    g671(.A(new_n530), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n532), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n534), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n532), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n682), .A4(new_n855), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT113), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n785), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(KEYINPUT114), .A3(new_n865), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n853), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n698), .B(new_n706), .C1(new_n705), .C2(new_n729), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n768), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n851), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n762), .B1(new_n722), .B2(new_n724), .ZN(new_n874));
  INV_X1    g688(.A(new_n869), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT114), .B1(new_n864), .B2(new_n865), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n768), .A4(new_n871), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(KEYINPUT116), .B(new_n827), .C1(new_n850), .C2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n755), .A2(new_n849), .A3(new_n838), .A4(new_n839), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n797), .A2(new_n833), .A3(new_n834), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n792), .A2(new_n793), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n789), .B1(new_n775), .B2(new_n776), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT52), .B1(new_n870), .B2(new_n872), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n879), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT53), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n879), .A3(new_n873), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT116), .B1(new_n892), .B2(new_n827), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n888), .A2(new_n879), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n827), .B1(new_n850), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n879), .A4(new_n873), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n725), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n778), .A2(new_n747), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n544), .A3(new_n328), .A4(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n656), .A3(new_n653), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n811), .A2(new_n328), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n905), .A2(new_n767), .A3(new_n902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n544), .A3(new_n760), .ZN(new_n907));
  INV_X1    g721(.A(new_n713), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n714), .B1(new_n909), .B2(KEYINPUT50), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n908), .A2(new_n747), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(KEYINPUT50), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n904), .B(new_n906), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n907), .A2(new_n778), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n734), .A2(new_n491), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n499), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n821), .A2(new_n822), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n912), .A2(new_n913), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n914), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n914), .A2(new_n921), .A3(KEYINPUT51), .A4(new_n922), .ZN(new_n926));
  OAI221_X1 g740(.A(new_n324), .B1(new_n903), .B2(new_n657), .C1(new_n907), .C2(new_n749), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n905), .A2(new_n777), .A3(new_n902), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT48), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(KEYINPUT48), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n900), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n916), .A2(KEYINPUT49), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n544), .A2(new_n337), .A3(new_n499), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n916), .A2(KEYINPUT49), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR4_X1    g751(.A1(new_n908), .A2(new_n809), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n933), .B1(new_n725), .B2(new_n938), .ZN(G75));
  NOR2_X1   g753(.A1(new_n253), .A2(G952), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n235), .B1(new_n896), .B2(new_n898), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT56), .B1(new_n942), .B2(G210), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n426), .A2(new_n429), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n427), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n941), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n943), .B2(new_n947), .ZN(G51));
  AND3_X1   g763(.A1(new_n942), .A2(new_n800), .A3(new_n802), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n486), .A2(new_n490), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT53), .B1(new_n887), .B2(new_n889), .ZN(new_n952));
  NOR4_X1   g766(.A1(new_n880), .A2(new_n882), .A3(new_n886), .A4(new_n827), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT54), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n899), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n492), .B(KEYINPUT57), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n950), .B1(new_n957), .B2(KEYINPUT119), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT119), .ZN(new_n959));
  INV_X1    g773(.A(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n954), .B2(new_n899), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(new_n951), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n940), .B1(new_n958), .B2(new_n962), .ZN(G54));
  NAND3_X1  g777(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .ZN(new_n964));
  INV_X1    g778(.A(new_n316), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n941), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT120), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G60));
  INV_X1    g783(.A(new_n955), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n242), .A2(new_n235), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(new_n974));
  OR2_X1    g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n941), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n900), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n971), .ZN(G63));
  NAND2_X1  g793(.A1(new_n896), .A2(new_n898), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n227), .A2(new_n235), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n681), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n940), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n980), .A2(new_n983), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n984), .B(new_n986), .C1(new_n987), .C2(new_n540), .ZN(new_n988));
  NAND2_X1  g802(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT124), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n988), .B(new_n991), .ZN(G66));
  INV_X1    g806(.A(new_n329), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n253), .B1(new_n993), .B2(G224), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n882), .B2(new_n253), .ZN(new_n995));
  INV_X1    g809(.A(G898), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n944), .B1(new_n996), .B2(G953), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G69));
  INV_X1    g812(.A(new_n872), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n726), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n625), .A2(new_n710), .A3(new_n778), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n847), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1002), .A2(new_n816), .A3(new_n825), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n253), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n305), .A2(new_n306), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n611), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n814), .A2(new_n815), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n777), .A2(new_n852), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n807), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n825), .A2(new_n795), .A3(new_n797), .A4(new_n999), .ZN(new_n1012));
  OR3_X1    g826(.A1(new_n1011), .A2(new_n1012), .A3(G953), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(G900), .B2(G953), .ZN(new_n1014));
  AOI22_X1  g828(.A1(new_n1006), .A2(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT125), .Z(new_n1017));
  XNOR2_X1  g831(.A(new_n1015), .B(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1005), .B2(new_n882), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n612), .A2(new_n578), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n588), .A2(new_n589), .A3(new_n607), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1011), .A2(new_n1012), .A3(new_n882), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1020), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1023), .A2(new_n941), .A3(new_n1027), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n891), .A2(new_n893), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT126), .Z(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1029), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1028), .B1(new_n1033), .B2(new_n1035), .ZN(G57));
endmodule


