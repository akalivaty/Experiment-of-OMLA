//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G250), .B1(G257), .B2(G264), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n208), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(new_n203), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT66), .B(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n203), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n222), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT67), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G50), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G50), .B2(new_n249), .ZN(new_n256));
  INV_X1    g0056(.A(new_n252), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n204), .A2(G20), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT8), .B(G58), .Z(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT68), .A2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT68), .A2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n267), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n215), .B1(KEYINPUT69), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G33), .A3(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(G226), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G222), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(G1698), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n287), .B1(new_n288), .B2(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n276), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT70), .B1(new_n293), .B2(new_n215), .ZN(new_n294));
  INV_X1    g0094(.A(new_n215), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(new_n276), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n273), .B(new_n281), .C1(new_n292), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n265), .B(new_n300), .C1(new_n301), .C2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(G190), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n265), .B(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n303), .B(new_n305), .C1(new_n306), .C2(new_n299), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n298), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n291), .A2(new_n223), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(G107), .B2(new_n285), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n286), .A2(G232), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n273), .B1(G244), .B2(new_n280), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G200), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n314), .B1(new_n319), .B2(new_n289), .C1(new_n223), .C2(new_n291), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n298), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G190), .A3(new_n316), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n257), .A2(new_n249), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n254), .A2(G77), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(G77), .B2(new_n249), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n259), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n327), .A2(KEYINPUT71), .B1(new_n261), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(KEYINPUT71), .B2(new_n327), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n326), .B1(new_n331), .B2(new_n252), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n318), .B(new_n322), .C1(new_n323), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n252), .ZN(new_n334));
  INV_X1    g0134(.A(new_n326), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n315), .B2(new_n317), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n321), .A2(new_n301), .A3(new_n316), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT73), .B1(new_n310), .B2(new_n344), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n280), .A2(G238), .B1(new_n269), .B2(new_n271), .ZN(new_n347));
  INV_X1    g0147(.A(G1698), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n282), .A2(new_n284), .A3(G226), .A4(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n282), .A2(new_n284), .A3(G232), .A4(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n298), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n347), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n347), .B2(new_n353), .ZN(new_n357));
  OAI21_X1  g0157(.A(G169), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(KEYINPUT75), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G169), .B(new_n360), .C1(new_n356), .C2(new_n357), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n353), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(G179), .A3(new_n355), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n366), .A2(new_n369), .A3(G179), .A4(new_n355), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n373));
  INV_X1    g0173(.A(G50), .ZN(new_n374));
  INV_X1    g0174(.A(new_n262), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n252), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT11), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT74), .B1(new_n249), .B2(G68), .ZN(new_n380));
  XOR2_X1   g0180(.A(new_n380), .B(KEYINPUT12), .Z(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n377), .B2(new_n378), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n372), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n366), .A2(G190), .A3(new_n355), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n356), .A2(new_n357), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n385), .B(new_n388), .C1(new_n389), .C2(new_n306), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n345), .A2(new_n346), .B1(KEYINPUT77), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n387), .ZN(new_n393));
  INV_X1    g0193(.A(new_n390), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT77), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  AOI21_X1  g0196(.A(G20), .B1(new_n282), .B2(new_n284), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT80), .B1(new_n397), .B2(KEYINPUT7), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT80), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n289), .C2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n284), .B1(new_n403), .B2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n400), .A2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n203), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G58), .A2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n217), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G20), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n262), .A2(G159), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n396), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n282), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n403), .B2(G33), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT7), .B1(new_n415), .B2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n283), .A2(KEYINPUT78), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n419), .A3(G33), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n282), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n400), .A3(new_n208), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n416), .A2(G68), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT79), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n410), .A2(new_n424), .A3(new_n411), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n208), .B1(new_n217), .B2(new_n408), .ZN(new_n426));
  INV_X1    g0226(.A(new_n411), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT79), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n425), .A2(new_n428), .A3(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n257), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n413), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n259), .A2(new_n254), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n432), .A2(new_n324), .B1(new_n249), .B2(new_n259), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT81), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n279), .A3(new_n295), .ZN(new_n438));
  INV_X1    g0238(.A(new_n275), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G232), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n272), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  MUX2_X1   g0243(.A(G223), .B(G226), .S(G1698), .Z(new_n444));
  NAND2_X1  g0244(.A1(new_n415), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G87), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n443), .B(G179), .C1(new_n447), .C2(new_n311), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n311), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g0249(.A(G169), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n435), .A2(new_n436), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G190), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n443), .B(new_n453), .C1(new_n447), .C2(new_n311), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n306), .B1(new_n449), .B2(new_n442), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n431), .A2(new_n434), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT81), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n433), .B(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n413), .B2(new_n430), .ZN(new_n462));
  INV_X1    g0262(.A(new_n451), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT18), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(KEYINPUT17), .A3(new_n456), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n452), .A2(new_n459), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n395), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n392), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT87), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G257), .A2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(G264), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(G1698), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n415), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n285), .A2(G303), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n311), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n274), .A2(new_n270), .A3(G1), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n438), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n207), .B(G45), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n438), .ZN(new_n484));
  INV_X1    g0284(.A(G270), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(G169), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n208), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G33), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT20), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n252), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT83), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n251), .A2(new_n215), .B1(G20), .B2(new_n493), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n488), .B(new_n208), .C1(G33), .C2(new_n490), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n252), .A3(new_n494), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n503), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n249), .A2(new_n493), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n257), .B(new_n249), .C1(G1), .C2(new_n260), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(new_n493), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n515), .A3(new_n512), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n487), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n471), .B1(new_n517), .B2(KEYINPUT21), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n508), .A2(new_n515), .A3(new_n512), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n515), .B1(new_n508), .B2(new_n512), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT87), .B(new_n519), .C1(new_n522), .C2(new_n487), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n477), .A2(new_n486), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G179), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n514), .B2(new_n516), .ZN(new_n527));
  OAI211_X1 g0327(.A(KEYINPUT21), .B(G169), .C1(new_n477), .C2(new_n486), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n520), .B2(new_n521), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT86), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(KEYINPUT86), .C1(new_n520), .C2(new_n521), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n525), .A2(G190), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n522), .B(new_n535), .C1(new_n306), .C2(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n524), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n249), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n511), .B2(G97), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(G97), .B(G107), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n490), .A3(G107), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n398), .A2(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n319), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n541), .B1(new_n550), .B2(new_n252), .ZN(new_n551));
  INV_X1    g0351(.A(G244), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G1698), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n420), .A2(new_n282), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(KEYINPUT4), .A2(G244), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n282), .A2(new_n284), .A3(new_n557), .A4(new_n348), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n558), .A2(new_n559), .A3(new_n488), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n311), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n483), .A2(new_n438), .A3(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n482), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n306), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n559), .A3(new_n488), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n555), .B2(new_n554), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n453), .C1(new_n567), .C2(new_n311), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n551), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n339), .B1(new_n561), .B2(new_n563), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n565), .B(new_n301), .C1(new_n567), .C2(new_n311), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n551), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n538), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n545), .B1(new_n543), .B2(new_n542), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n208), .B1(new_n288), .B2(new_n375), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n402), .A2(new_n406), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n540), .B1(new_n579), .B2(new_n257), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n572), .A3(new_n571), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n551), .A2(new_n569), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(KEYINPUT82), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n415), .A2(KEYINPUT88), .A3(new_n208), .A4(G87), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n420), .A2(new_n208), .A3(G87), .A4(new_n282), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  OR4_X1    g0390(.A1(KEYINPUT22), .A2(new_n285), .A3(G20), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n208), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n319), .A2(KEYINPUT23), .A3(G20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n594), .A2(new_n595), .B1(new_n597), .B2(new_n208), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT24), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n257), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT25), .B1(new_n250), .B2(new_n319), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n511), .A2(G107), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  MUX2_X1   g0409(.A(G250), .B(G257), .S(G1698), .Z(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n420), .A3(new_n282), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G294), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n297), .B2(new_n294), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n484), .A2(new_n473), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n482), .ZN(new_n616));
  INV_X1    g0416(.A(new_n482), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n613), .A2(new_n614), .A3(new_n617), .A4(KEYINPUT89), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n616), .A2(new_n339), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n482), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n301), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n603), .A2(new_n608), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n602), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n601), .B1(new_n592), .B2(new_n598), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n252), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n453), .B1(new_n616), .B2(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n306), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n628), .A3(new_n607), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT19), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n261), .A2(new_n630), .A3(G97), .ZN(new_n631));
  NOR2_X1   g0431(.A1(G97), .A2(G107), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n590), .B1(new_n351), .B2(new_n208), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n630), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n420), .A2(new_n208), .A3(G68), .A4(new_n282), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n252), .B1(new_n250), .B2(new_n328), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n511), .A2(new_n329), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(G238), .A2(G1698), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n552), .B2(G1698), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n420), .A3(new_n282), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n596), .B1(new_n297), .B2(new_n294), .ZN(new_n643));
  INV_X1    g0443(.A(new_n481), .ZN(new_n644));
  OAI21_X1  g0444(.A(G250), .B1(new_n274), .B2(G1), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n438), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n339), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n438), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n597), .B1(new_n415), .B2(new_n641), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n301), .B(new_n649), .C1(new_n650), .C2(new_n311), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n639), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(G200), .B1(new_n643), .B2(new_n647), .ZN(new_n653));
  OAI211_X1 g0453(.A(G190), .B(new_n649), .C1(new_n650), .C2(new_n311), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n511), .A2(G87), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n637), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n584), .A2(new_n622), .A3(new_n629), .A4(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n470), .A2(new_n537), .A3(new_n659), .ZN(G372));
  AOI21_X1  g0460(.A(new_n393), .B1(new_n390), .B2(new_n343), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n459), .A2(new_n465), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n464), .B(new_n452), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n308), .A2(new_n309), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n302), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT93), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT92), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n580), .A2(new_n667), .A3(new_n572), .A4(new_n571), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT92), .B1(new_n551), .B2(new_n573), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n648), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n649), .B1(new_n650), .B2(new_n311), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n339), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n651), .A3(new_n639), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n668), .A2(new_n669), .A3(new_n675), .A4(new_n656), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n675), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n657), .A2(new_n551), .A3(new_n573), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n524), .A2(new_n534), .A3(new_n622), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n581), .A2(new_n675), .A3(new_n656), .A4(new_n582), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n603), .A2(new_n608), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n628), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n682), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n666), .B1(new_n470), .B2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G343), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT94), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n522), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n537), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n524), .A2(new_n534), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n622), .A2(new_n629), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n685), .B2(new_n699), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n622), .A2(new_n699), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n622), .A2(new_n698), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n698), .B1(new_n524), .B2(new_n534), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(G399));
  NOR2_X1   g0515(.A1(new_n212), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR4_X1   g0517(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n218), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n691), .B2(new_n698), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT96), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT26), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n678), .B1(new_n679), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n683), .B2(new_n686), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n725), .B1(new_n730), .B2(new_n698), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n726), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n687), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT96), .A3(new_n699), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g0536(.A(new_n682), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n683), .A2(new_n689), .A3(new_n686), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n689), .B1(new_n683), .B2(new_n686), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n699), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n722), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n724), .A2(new_n736), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n524), .A2(new_n534), .A3(new_n536), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n657), .B1(new_n575), .B2(new_n583), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n706), .A3(new_n746), .A4(new_n699), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n643), .A2(new_n647), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n525), .A2(G179), .A3(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n749), .B(new_n620), .C1(new_n561), .C2(new_n563), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n561), .A2(new_n563), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n615), .A3(new_n748), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n753), .B2(new_n526), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n753), .A2(new_n526), .A3(new_n751), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n698), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n744), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n721), .B1(new_n762), .B2(G1), .ZN(G364));
  AND2_X1   g0563(.A1(new_n208), .A2(G13), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n207), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n716), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n705), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n704), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n215), .B1(G20), .B2(new_n339), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n208), .A2(new_n301), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  NAND3_X1  g0577(.A1(new_n773), .A2(G190), .A3(new_n306), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT101), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n208), .A2(G179), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT99), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n782), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT100), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G329), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n782), .A2(new_n453), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(new_n790), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n453), .A2(G179), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n208), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n285), .B1(new_n797), .B2(new_n798), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n774), .A2(new_n453), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n796), .B(new_n802), .C1(G326), .C2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n781), .A2(new_n789), .A3(new_n793), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n794), .A2(new_n319), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n289), .B1(new_n797), .B2(new_n288), .C1(new_n202), .C2(new_n778), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G68), .C2(new_n775), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n788), .A2(G87), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n791), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n813));
  INV_X1    g0613(.A(new_n800), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(G97), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n803), .A2(G50), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n808), .A2(new_n809), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n772), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n771), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n211), .A2(new_n289), .ZN(new_n824));
  INV_X1    g0624(.A(G355), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n825), .B1(G116), .B2(new_n211), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT97), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n247), .A2(new_n274), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n212), .A2(new_n415), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n266), .A2(new_n268), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n219), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n827), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n770), .B(new_n819), .C1(new_n823), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n822), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n704), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n769), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n342), .A2(new_n698), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n332), .B2(new_n699), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n336), .A2(KEYINPUT104), .A3(new_n698), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n337), .C2(new_n333), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n843), .B2(new_n342), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n741), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n698), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n740), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n767), .B1(new_n849), .B2(new_n760), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n760), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n771), .A2(new_n820), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n770), .B1(new_n288), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n794), .A2(new_n590), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n792), .B2(G311), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n800), .A2(new_n490), .B1(new_n778), .B2(new_n801), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT103), .ZN(new_n858));
  INV_X1    g0658(.A(new_n797), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n289), .B1(new_n859), .B2(G116), .ZN(new_n860));
  INV_X1    g0660(.A(new_n803), .ZN(new_n861));
  INV_X1    g0661(.A(G303), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .C1(new_n795), .C2(new_n776), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n858), .B(new_n863), .C1(G107), .C2(new_n788), .ZN(new_n864));
  INV_X1    g0664(.A(new_n778), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(G143), .B1(new_n859), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n861), .B2(new_n867), .C1(new_n868), .C2(new_n776), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n415), .B1(new_n203), .B2(new_n794), .C1(new_n202), .C2(new_n800), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n787), .A2(new_n374), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(G132), .C2(new_n792), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n856), .A2(new_n864), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n853), .B1(new_n772), .B2(new_n874), .C1(new_n844), .C2(new_n821), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n851), .A2(new_n876), .ZN(G384));
  OR2_X1    g0677(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n216), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  NAND3_X1  g0681(.A1(new_n219), .A2(G77), .A3(new_n408), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n201), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n207), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n452), .A2(new_n464), .ZN(new_n886));
  INV_X1    g0686(.A(new_n696), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n423), .A2(new_n429), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n252), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n425), .A2(new_n428), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n423), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n434), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n451), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n696), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n457), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n435), .A2(KEYINPUT107), .A3(new_n451), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT107), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n462), .B2(new_n463), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n435), .A2(new_n696), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT37), .B1(new_n462), .B2(new_n456), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n895), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n466), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n457), .B(KEYINPUT108), .C1(new_n462), .C2(new_n463), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n901), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n435), .A2(new_n451), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT108), .B1(new_n915), .B2(new_n457), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n901), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n917), .A2(new_n903), .B1(new_n466), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n912), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n911), .B1(new_n921), .B2(KEYINPUT39), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n387), .A2(new_n698), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n888), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n839), .ZN(new_n926));
  INV_X1    g0726(.A(new_n847), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n691), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n364), .A2(new_n371), .A3(new_n390), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n699), .A2(new_n385), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n931), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n362), .A2(new_n363), .B1(new_n368), .B2(new_n370), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n390), .B(new_n933), .C1(new_n934), .C2(new_n385), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n387), .A2(new_n929), .A3(new_n390), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n907), .A2(new_n908), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n925), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n724), .A2(new_n469), .A3(new_n736), .A4(new_n743), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n666), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n943), .B(new_n945), .Z(new_n946));
  AND2_X1   g0746(.A1(new_n469), .A2(new_n759), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n936), .A2(new_n844), .A3(new_n937), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n659), .A2(new_n537), .A3(new_n698), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT31), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n757), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n948), .B1(new_n953), .B2(new_n941), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n936), .A2(new_n844), .A3(new_n937), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n747), .B2(new_n758), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n920), .A2(new_n956), .A3(KEYINPUT40), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n947), .A2(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(G330), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n207), .B2(new_n764), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n946), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n885), .B1(new_n963), .B2(new_n964), .ZN(G367));
  OAI211_X1 g0765(.A(new_n581), .B(new_n582), .C1(new_n551), .C2(new_n699), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n574), .A2(new_n698), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n713), .A2(new_n706), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n581), .B1(new_n967), .B2(new_n622), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n699), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n637), .A2(new_n655), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n698), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n675), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n675), .A2(new_n656), .A3(new_n977), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n972), .A2(new_n984), .A3(new_n974), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n983), .B2(new_n985), .ZN(new_n987));
  INV_X1    g0787(.A(new_n969), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n705), .A2(new_n710), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n987), .B1(KEYINPUT111), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n970), .B1(new_n710), .B2(new_n713), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n705), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n997), .A2(new_n761), .A3(KEYINPUT112), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT112), .B1(new_n997), .B2(new_n761), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n988), .A2(new_n714), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n714), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n969), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT45), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1001), .A2(new_n711), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n711), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n998), .A2(new_n999), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT113), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n998), .A2(KEYINPUT113), .A3(new_n999), .A4(new_n1007), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n761), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n716), .B(KEYINPUT41), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n765), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n994), .A2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n800), .A2(new_n203), .B1(new_n794), .B2(new_n288), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n289), .B1(new_n791), .B2(new_n867), .C1(new_n778), .C2(new_n868), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(G143), .C2(new_n803), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n201), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n775), .A2(G159), .B1(new_n859), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT115), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(new_n202), .C2(new_n787), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n788), .A2(G116), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT46), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT114), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n861), .A2(new_n798), .B1(new_n319), .B2(new_n800), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n415), .B1(new_n775), .B2(G294), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n791), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n865), .A2(G303), .B1(new_n1030), .B2(G317), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n795), .C2(new_n797), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n794), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1028), .B(new_n1032), .C1(G97), .C2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1023), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT47), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n771), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n978), .A2(new_n822), .A3(new_n979), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n829), .A2(new_n240), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n823), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n212), .B2(new_n329), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n770), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1015), .A2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n998), .A2(new_n999), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n717), .B1(new_n997), .B2(new_n761), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n709), .A2(new_n822), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n237), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n829), .B1(new_n1050), .B2(new_n830), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n718), .B2(new_n824), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n259), .A2(new_n374), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT50), .Z(new_n1054));
  AOI21_X1  g0854(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n718), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1052), .A2(new_n1056), .B1(new_n319), .B2(new_n212), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n767), .B1(new_n1057), .B2(new_n1041), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n800), .A2(new_n328), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n810), .B2(new_n861), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n259), .B2(new_n775), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n797), .A2(new_n203), .B1(new_n791), .B2(new_n868), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n415), .B1(new_n490), .B2(new_n794), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G50), .C2(new_n865), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n788), .A2(G77), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n415), .B1(G326), .B2(new_n1030), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n801), .B1(new_n795), .B2(new_n800), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n865), .A2(G317), .B1(new_n859), .B2(G303), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n861), .B2(new_n779), .C1(new_n798), .C2(new_n776), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1068), .B1(new_n493), .B2(new_n794), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT117), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n772), .B1(new_n1078), .B2(KEYINPUT117), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1058), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n996), .A2(new_n766), .B1(new_n1049), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1048), .A2(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(G393));
  INV_X1    g0886(.A(new_n829), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n823), .B1(new_n490), .B2(new_n211), .C1(new_n1087), .C2(new_n244), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n767), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n806), .B1(G116), .B2(new_n814), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n862), .B2(new_n776), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n787), .A2(new_n795), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n285), .B1(new_n791), .B2(new_n779), .C1(new_n797), .C2(new_n801), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G317), .A2(new_n803), .B1(new_n865), .B2(G311), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n800), .A2(new_n288), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n854), .B(new_n1097), .C1(new_n1019), .C2(new_n775), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n788), .A2(G68), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n259), .A2(new_n859), .B1(new_n1030), .B2(G143), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n415), .A4(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G150), .A2(new_n803), .B1(new_n865), .B2(G159), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1094), .A2(new_n1096), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n1104), .B2(new_n771), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n988), .B2(new_n835), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1007), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n765), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n717), .B1(new_n1046), .B2(new_n1107), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  OAI21_X1  g0912(.A(new_n938), .B1(new_n760), .B2(new_n845), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n759), .A2(G330), .A3(new_n844), .A4(new_n939), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(new_n926), .B2(new_n848), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n843), .A2(new_n342), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n839), .B1(new_n735), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n469), .A2(G330), .A3(new_n759), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n944), .A2(new_n666), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n920), .A2(new_n924), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT96), .B1(new_n733), .B2(new_n699), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n725), .B(new_n698), .C1(new_n687), .C2(new_n732), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1116), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n926), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1129), .B2(new_n939), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n910), .B1(new_n909), .B2(new_n920), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n940), .B2(new_n924), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1124), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1117), .B2(new_n938), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n938), .B1(new_n848), .B2(new_n926), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n922), .B1(new_n1136), .B2(new_n923), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1137), .A3(new_n1114), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1123), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1135), .A2(new_n1137), .A3(new_n1114), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1114), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1122), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1144), .A3(new_n716), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1133), .A2(new_n766), .A3(new_n1138), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT119), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT119), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1133), .A2(new_n1148), .A3(new_n766), .A4(new_n1138), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n776), .A2(new_n319), .B1(new_n861), .B2(new_n795), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1097), .B(new_n1151), .C1(G68), .C2(new_n1033), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n792), .A2(G294), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n285), .B1(new_n778), .B2(new_n493), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G97), .B2(new_n859), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1152), .A2(new_n809), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n776), .A2(new_n867), .B1(new_n861), .B2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n800), .A2(new_n810), .B1(new_n794), .B2(new_n201), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT53), .B1(new_n787), .B2(new_n868), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n792), .A2(G125), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n797), .A2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n285), .B(new_n1164), .C1(G132), .C2(new_n865), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n868), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1156), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n771), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n259), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n770), .B1(new_n1170), .B2(new_n852), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n1131), .C2(new_n821), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT120), .B1(new_n1150), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1172), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1145), .B1(new_n1173), .B2(new_n1176), .ZN(G378));
  NAND3_X1  g0977(.A1(new_n954), .A2(new_n957), .A3(G330), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT124), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT123), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n310), .B(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n265), .A2(new_n887), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT55), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1184), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1183), .B(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1180), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1183), .B(new_n1187), .Z(new_n1190));
  NAND4_X1  g0990(.A1(new_n958), .A2(new_n1190), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n943), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1189), .A2(new_n943), .A3(new_n1191), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n766), .A3(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n861), .A2(new_n493), .B1(new_n203), .B2(new_n800), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT121), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n794), .A2(new_n202), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n778), .A2(new_n319), .B1(new_n797), .B2(new_n328), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G97), .C2(new_n775), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G41), .B(new_n415), .C1(new_n792), .C2(G283), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1201), .A3(new_n1066), .A4(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT58), .Z(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n260), .B2(new_n267), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n415), .B2(G41), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n778), .A2(new_n1157), .B1(new_n797), .B2(new_n867), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G132), .B2(new_n775), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G150), .A2(new_n814), .B1(new_n803), .B2(G125), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n787), .C2(new_n1163), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1033), .A2(G159), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n1030), .C2(G124), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1206), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n771), .B1(new_n1204), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n770), .B1(new_n201), .B2(new_n852), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n1188), .C2(new_n821), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1196), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1121), .B1(new_n1143), .B2(new_n1122), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n716), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1195), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n943), .B1(new_n1191), .B2(new_n1189), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1121), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1139), .B2(new_n1119), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1221), .B1(new_n1224), .B2(new_n1230), .ZN(G375));
  OR2_X1    g1031(.A1(new_n1119), .A2(new_n765), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G116), .A2(new_n775), .B1(new_n803), .B2(G294), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n1060), .C1(new_n288), .C2(new_n794), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n289), .B1(new_n859), .B2(G107), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n792), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1235), .B1(new_n795), .B2(new_n778), .C1(new_n1236), .C2(new_n862), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(G97), .C2(new_n788), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1199), .B1(G50), .B2(new_n814), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n803), .A2(G132), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n776), .C2(new_n1163), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n865), .A2(G137), .B1(new_n859), .B2(G150), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n415), .C1(new_n1236), .C2(new_n1157), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(G159), .C2(new_n788), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n771), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n770), .B1(new_n203), .B2(new_n852), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n939), .C2(new_n821), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1232), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1013), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1123), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G381));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OR3_X1    g1054(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1255));
  OR2_X1    g1055(.A1(G378), .A2(G375), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G387), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1058(.A1(G378), .A2(G375), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1222), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1220), .B1(new_n1261), .B2(new_n1249), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1145), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1250), .B1(new_n1122), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1119), .A2(new_n1121), .A3(KEYINPUT60), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n716), .A3(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1270), .A2(G384), .A3(new_n1248), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1270), .B2(new_n1248), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1259), .A2(new_n1263), .A3(new_n1266), .A4(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1145), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1150), .A2(new_n1172), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1174), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n1172), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1265), .B1(new_n1281), .B2(new_n1262), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1275), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1282), .A2(new_n1273), .A3(new_n1259), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1276), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1265), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1259), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1273), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1293), .A3(new_n1289), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT125), .B1(new_n1273), .B2(new_n1288), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1287), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT127), .B1(new_n1286), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1273), .B1(new_n1282), .B2(new_n1259), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1295), .B(new_n1294), .C1(new_n1299), .C2(new_n1289), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1276), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .A4(new_n1287), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G390), .B1(new_n1015), .B2(new_n1044), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1044), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1305), .B(new_n1111), .C1(new_n994), .C2(new_n1014), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n837), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n1304), .A2(new_n1306), .B1(new_n1253), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(new_n1111), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1253), .A2(new_n1307), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1015), .A2(new_n1044), .A3(G390), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1298), .A2(new_n1303), .A3(new_n1313), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1274), .B(KEYINPUT63), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1315), .A2(new_n1287), .A3(new_n1300), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1291), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1313), .B(new_n1320), .ZN(G402));
endmodule


