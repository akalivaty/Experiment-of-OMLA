

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U554 ( .A1(n639), .A2(n913), .ZN(n638) );
  INV_X1 U555 ( .A(G2104), .ZN(n531) );
  OR2_X1 U556 ( .A1(n715), .A2(n714), .ZN(n523) );
  BUF_X1 U557 ( .A(n896), .Z(n524) );
  NOR2_X1 U558 ( .A1(G2105), .A2(n531), .ZN(n896) );
  BUF_X2 U559 ( .A(n897), .Z(n525) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n534), .Z(n897) );
  NOR2_X1 U561 ( .A1(n622), .A2(n992), .ZN(n624) );
  AND2_X1 U562 ( .A1(n653), .A2(G1996), .ZN(n609) );
  BUF_X1 U563 ( .A(n658), .Z(n678) );
  INV_X1 U564 ( .A(n658), .ZN(n653) );
  NAND2_X1 U565 ( .A1(n607), .A2(n716), .ZN(n658) );
  NOR2_X2 U566 ( .A1(n531), .A2(n535), .ZN(n900) );
  XNOR2_X1 U567 ( .A(n659), .B(KEYINPUT97), .ZN(n713) );
  NOR2_X1 U568 ( .A1(n619), .A2(n618), .ZN(n621) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n529) );
  NOR2_X1 U570 ( .A1(n747), .A2(n755), .ZN(n526) );
  XOR2_X1 U571 ( .A(KEYINPUT102), .B(n672), .Z(n527) );
  NOR2_X1 U572 ( .A1(n693), .A2(n692), .ZN(n528) );
  INV_X1 U573 ( .A(KEYINPUT26), .ZN(n608) );
  INV_X1 U574 ( .A(G8), .ZN(n660) );
  OR2_X1 U575 ( .A1(n673), .A2(n660), .ZN(n661) );
  NOR2_X1 U576 ( .A1(n667), .A2(n666), .ZN(n668) );
  INV_X1 U577 ( .A(KEYINPUT32), .ZN(n685) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  NOR2_X1 U579 ( .A1(G651), .A2(n580), .ZN(n801) );
  XNOR2_X1 U580 ( .A(n530), .B(n529), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G101), .A2(n896), .ZN(n530) );
  INV_X1 U582 ( .A(G2105), .ZN(n535) );
  NAND2_X1 U583 ( .A1(n900), .A2(G113), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U585 ( .A1(G137), .A2(n525), .ZN(n537) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n535), .ZN(n901) );
  NAND2_X1 U587 ( .A1(G125), .A2(n901), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U589 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n807) );
  NAND2_X1 U591 ( .A1(G91), .A2(n807), .ZN(n541) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n580) );
  XNOR2_X1 U593 ( .A(KEYINPUT65), .B(G651), .ZN(n545) );
  NOR2_X1 U594 ( .A1(n580), .A2(n545), .ZN(n808) );
  NAND2_X1 U595 ( .A1(G78), .A2(n808), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n801), .A2(G53), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT70), .B(n542), .Z(n543) );
  NOR2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NOR2_X1 U600 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X2 U601 ( .A(KEYINPUT1), .B(n546), .Z(n803) );
  NAND2_X1 U602 ( .A1(G65), .A2(n803), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U604 ( .A1(G90), .A2(n807), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G77), .A2(n808), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(KEYINPUT9), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n552), .B(n551), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n801), .A2(G52), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G64), .A2(n803), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(KEYINPUT68), .B(n555), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U614 ( .A(G171), .ZN(G301) );
  NAND2_X1 U615 ( .A1(n801), .A2(G51), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G63), .A2(n803), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U618 ( .A(KEYINPUT6), .B(n560), .ZN(n567) );
  NAND2_X1 U619 ( .A1(n807), .A2(G89), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G76), .A2(n808), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n564), .ZN(n565) );
  XNOR2_X1 U624 ( .A(KEYINPUT77), .B(n565), .ZN(n566) );
  NOR2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(n568), .Z(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(n808), .A2(G75), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT86), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n801), .A2(G50), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G62), .A2(n803), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G88), .A2(n807), .ZN(n572) );
  XNOR2_X1 U634 ( .A(KEYINPUT85), .B(n572), .ZN(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G303) );
  INV_X1 U637 ( .A(G303), .ZN(G166) );
  NAND2_X1 U638 ( .A1(G49), .A2(n801), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U641 ( .A(n579), .B(KEYINPUT83), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G87), .A2(n580), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n803), .A2(n583), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT84), .B(n584), .Z(G288) );
  NAND2_X1 U646 ( .A1(n807), .A2(G86), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G61), .A2(n803), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n808), .A2(G73), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n801), .A2(G48), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G72), .A2(n808), .ZN(n598) );
  NAND2_X1 U655 ( .A1(G85), .A2(n807), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G47), .A2(n801), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U658 ( .A1(n803), .A2(G60), .ZN(n594) );
  XOR2_X1 U659 ( .A(KEYINPUT66), .B(n594), .Z(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U662 ( .A(KEYINPUT67), .B(n599), .Z(G290) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n717) );
  INV_X1 U664 ( .A(n717), .ZN(n607) );
  NAND2_X1 U665 ( .A1(n900), .A2(G114), .ZN(n600) );
  XNOR2_X1 U666 ( .A(n600), .B(KEYINPUT92), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G102), .A2(n524), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U669 ( .A1(G126), .A2(n901), .ZN(n604) );
  NAND2_X1 U670 ( .A1(G138), .A2(n525), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U672 ( .A1(n606), .A2(n605), .ZN(n773) );
  NOR2_X2 U673 ( .A1(n773), .A2(G1384), .ZN(n716) );
  XNOR2_X1 U674 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U675 ( .A1(n678), .A2(G1341), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n611), .A2(n610), .ZN(n622) );
  XNOR2_X1 U677 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n616) );
  NAND2_X1 U678 ( .A1(n807), .A2(G81), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U680 ( .A1(G68), .A2(n808), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U682 ( .A(n616), .B(n615), .ZN(n619) );
  NAND2_X1 U683 ( .A1(G56), .A2(n803), .ZN(n617) );
  XOR2_X1 U684 ( .A(KEYINPUT14), .B(n617), .Z(n618) );
  NAND2_X1 U685 ( .A1(n801), .A2(G43), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n621), .A2(n620), .ZN(n992) );
  INV_X1 U687 ( .A(KEYINPUT64), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n624), .B(n623), .ZN(n639) );
  NAND2_X1 U689 ( .A1(G54), .A2(n801), .ZN(n631) );
  NAND2_X1 U690 ( .A1(G66), .A2(n803), .ZN(n626) );
  NAND2_X1 U691 ( .A1(G79), .A2(n808), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U693 ( .A1(G92), .A2(n807), .ZN(n627) );
  XNOR2_X1 U694 ( .A(KEYINPUT75), .B(n627), .ZN(n628) );
  NOR2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U697 ( .A(n632), .B(KEYINPUT15), .ZN(n633) );
  XNOR2_X1 U698 ( .A(KEYINPUT76), .B(n633), .ZN(n985) );
  INV_X1 U699 ( .A(n985), .ZN(n913) );
  NAND2_X1 U700 ( .A1(G1348), .A2(n678), .ZN(n635) );
  NAND2_X1 U701 ( .A1(G2067), .A2(n653), .ZN(n634) );
  NAND2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U703 ( .A(n636), .B(KEYINPUT100), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U705 ( .A1(n913), .A2(n639), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n646) );
  INV_X1 U707 ( .A(G299), .ZN(n979) );
  NAND2_X1 U708 ( .A1(n653), .A2(G2072), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT27), .ZN(n644) );
  AND2_X1 U710 ( .A1(G1956), .A2(n678), .ZN(n643) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U712 ( .A1(n979), .A2(n647), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n651) );
  NOR2_X1 U714 ( .A1(n979), .A2(n647), .ZN(n649) );
  XNOR2_X1 U715 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT29), .ZN(n657) );
  XOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .Z(n1006) );
  NOR2_X1 U720 ( .A1(n1006), .A2(n678), .ZN(n655) );
  NOR2_X1 U721 ( .A1(n653), .A2(G1961), .ZN(n654) );
  NOR2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n665) );
  NOR2_X1 U723 ( .A1(G301), .A2(n665), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n670) );
  XNOR2_X1 U725 ( .A(KEYINPUT101), .B(KEYINPUT30), .ZN(n663) );
  NAND2_X1 U726 ( .A1(n658), .A2(G8), .ZN(n659) );
  INV_X1 U727 ( .A(n713), .ZN(n693) );
  NOR2_X1 U728 ( .A1(G1966), .A2(n693), .ZN(n671) );
  NOR2_X1 U729 ( .A1(G2084), .A2(n678), .ZN(n673) );
  OR2_X1 U730 ( .A1(n671), .A2(n661), .ZN(n662) );
  XOR2_X1 U731 ( .A(n663), .B(n662), .Z(n664) );
  NOR2_X1 U732 ( .A1(G168), .A2(n664), .ZN(n667) );
  AND2_X1 U733 ( .A1(G301), .A2(n665), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n668), .B(KEYINPUT31), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n675), .A2(n671), .ZN(n672) );
  AND2_X1 U737 ( .A1(G8), .A2(n673), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n527), .A2(n674), .ZN(n688) );
  INV_X1 U739 ( .A(n675), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(G286), .ZN(n683) );
  NOR2_X1 U741 ( .A1(G1971), .A2(n693), .ZN(n677) );
  XNOR2_X1 U742 ( .A(KEYINPUT103), .B(n677), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n678), .ZN(n679) );
  NOR2_X1 U744 ( .A1(G166), .A2(n679), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n684), .A2(G8), .ZN(n686) );
  XNOR2_X1 U748 ( .A(n686), .B(n685), .ZN(n687) );
  OR2_X2 U749 ( .A1(n688), .A2(n687), .ZN(n708) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NOR2_X1 U752 ( .A1(n689), .A2(n984), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n708), .A2(n690), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n691), .B(KEYINPUT104), .ZN(n694) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U756 ( .A(n980), .ZN(n692) );
  AND2_X1 U757 ( .A1(n694), .A2(n528), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n695), .A2(KEYINPUT33), .ZN(n696) );
  XNOR2_X1 U759 ( .A(n696), .B(KEYINPUT105), .ZN(n702) );
  OR2_X1 U760 ( .A1(G1981), .A2(G305), .ZN(n703) );
  NAND2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n703), .A2(n697), .ZN(n996) );
  INV_X1 U763 ( .A(n996), .ZN(n700) );
  AND2_X1 U764 ( .A1(KEYINPUT33), .A2(n984), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n698), .A2(n713), .ZN(n699) );
  AND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n707) );
  XOR2_X1 U768 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT98), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n705), .A2(n713), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n715) );
  INV_X1 U772 ( .A(n708), .ZN(n711) );
  NAND2_X1 U773 ( .A1(G166), .A2(G8), .ZN(n709) );
  NOR2_X1 U774 ( .A1(G2090), .A2(n709), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(KEYINPUT93), .ZN(n758) );
  XNOR2_X1 U779 ( .A(G1986), .B(G290), .ZN(n983) );
  NAND2_X1 U780 ( .A1(G95), .A2(n524), .ZN(n720) );
  NAND2_X1 U781 ( .A1(G131), .A2(n525), .ZN(n719) );
  NAND2_X1 U782 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n900), .A2(G107), .ZN(n721) );
  XOR2_X1 U784 ( .A(KEYINPUT96), .B(n721), .Z(n722) );
  NOR2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U786 ( .A1(n901), .A2(G119), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n725), .A2(n724), .ZN(n893) );
  NAND2_X1 U788 ( .A1(G1991), .A2(n893), .ZN(n734) );
  NAND2_X1 U789 ( .A1(G117), .A2(n900), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G141), .A2(n525), .ZN(n726) );
  NAND2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U792 ( .A1(n524), .A2(G105), .ZN(n728) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(n728), .Z(n729) );
  NOR2_X1 U794 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U795 ( .A1(n901), .A2(G129), .ZN(n731) );
  NAND2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n877) );
  NAND2_X1 U797 ( .A1(G1996), .A2(n877), .ZN(n733) );
  NAND2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n961) );
  NOR2_X1 U799 ( .A1(n983), .A2(n961), .ZN(n735) );
  NOR2_X1 U800 ( .A1(n758), .A2(n735), .ZN(n747) );
  NAND2_X1 U801 ( .A1(G116), .A2(n900), .ZN(n737) );
  NAND2_X1 U802 ( .A1(G128), .A2(n901), .ZN(n736) );
  NAND2_X1 U803 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U804 ( .A(n738), .B(KEYINPUT35), .ZN(n744) );
  XNOR2_X1 U805 ( .A(KEYINPUT95), .B(KEYINPUT34), .ZN(n742) );
  NAND2_X1 U806 ( .A1(G104), .A2(n524), .ZN(n740) );
  NAND2_X1 U807 ( .A1(G140), .A2(n525), .ZN(n739) );
  NAND2_X1 U808 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U809 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U811 ( .A(KEYINPUT36), .B(n745), .ZN(n909) );
  XOR2_X1 U812 ( .A(G2067), .B(KEYINPUT37), .Z(n746) );
  XNOR2_X1 U813 ( .A(KEYINPUT94), .B(n746), .ZN(n748) );
  NAND2_X1 U814 ( .A1(n909), .A2(n748), .ZN(n968) );
  NOR2_X1 U815 ( .A1(n968), .A2(n758), .ZN(n755) );
  NAND2_X1 U816 ( .A1(n523), .A2(n526), .ZN(n761) );
  NOR2_X1 U817 ( .A1(n909), .A2(n748), .ZN(n957) );
  NOR2_X1 U818 ( .A1(n877), .A2(G1996), .ZN(n749) );
  XNOR2_X1 U819 ( .A(n749), .B(KEYINPUT106), .ZN(n952) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n893), .ZN(n955) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U822 ( .A1(n955), .A2(n750), .ZN(n751) );
  NOR2_X1 U823 ( .A1(n961), .A2(n751), .ZN(n752) );
  NOR2_X1 U824 ( .A1(n952), .A2(n752), .ZN(n753) );
  XOR2_X1 U825 ( .A(KEYINPUT39), .B(n753), .Z(n754) );
  NOR2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U827 ( .A1(n957), .A2(n756), .ZN(n757) );
  NOR2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U829 ( .A(n759), .B(KEYINPUT107), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U831 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U832 ( .A(G2451), .B(G2454), .Z(n764) );
  XNOR2_X1 U833 ( .A(G2430), .B(KEYINPUT108), .ZN(n763) );
  XNOR2_X1 U834 ( .A(n764), .B(n763), .ZN(n765) );
  XOR2_X1 U835 ( .A(n765), .B(G2446), .Z(n767) );
  XNOR2_X1 U836 ( .A(G1341), .B(G1348), .ZN(n766) );
  XNOR2_X1 U837 ( .A(n767), .B(n766), .ZN(n771) );
  XOR2_X1 U838 ( .A(G2438), .B(G2427), .Z(n769) );
  XNOR2_X1 U839 ( .A(G2443), .B(G2435), .ZN(n768) );
  XNOR2_X1 U840 ( .A(n769), .B(n768), .ZN(n770) );
  XOR2_X1 U841 ( .A(n771), .B(n770), .Z(n772) );
  AND2_X1 U842 ( .A1(G14), .A2(n772), .ZN(G401) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U844 ( .A(n773), .Z(G164) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  INV_X1 U848 ( .A(G108), .ZN(G238) );
  INV_X1 U849 ( .A(G120), .ZN(G236) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U851 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n776) );
  XNOR2_X1 U853 ( .A(G223), .B(KEYINPUT71), .ZN(n842) );
  NAND2_X1 U854 ( .A1(G567), .A2(n842), .ZN(n775) );
  XNOR2_X1 U855 ( .A(n776), .B(n775), .ZN(G234) );
  INV_X1 U856 ( .A(G860), .ZN(n782) );
  OR2_X1 U857 ( .A1(n992), .A2(n782), .ZN(G153) );
  NAND2_X1 U858 ( .A1(G301), .A2(G868), .ZN(n777) );
  XNOR2_X1 U859 ( .A(n777), .B(KEYINPUT74), .ZN(n779) );
  INV_X1 U860 ( .A(G868), .ZN(n823) );
  NAND2_X1 U861 ( .A1(n823), .A2(n913), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(G284) );
  NOR2_X1 U863 ( .A1(G286), .A2(n823), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G297) );
  NAND2_X1 U866 ( .A1(n782), .A2(G559), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n783), .A2(n985), .ZN(n784) );
  XNOR2_X1 U868 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(n913), .A2(n823), .ZN(n785) );
  XOR2_X1 U870 ( .A(KEYINPUT78), .B(n785), .Z(n786) );
  NOR2_X1 U871 ( .A1(G559), .A2(n786), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G868), .A2(n992), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G111), .A2(n900), .ZN(n790) );
  NAND2_X1 U875 ( .A1(G99), .A2(n524), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n797) );
  NAND2_X1 U877 ( .A1(G135), .A2(n525), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT80), .ZN(n795) );
  XOR2_X1 U879 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n793) );
  NAND2_X1 U880 ( .A1(G123), .A2(n901), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n793), .B(n792), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n954) );
  XNOR2_X1 U884 ( .A(n954), .B(G2096), .ZN(n799) );
  INV_X1 U885 ( .A(G2100), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(G156) );
  NAND2_X1 U887 ( .A1(n985), .A2(G559), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n800), .B(n992), .ZN(n820) );
  NOR2_X1 U889 ( .A1(n820), .A2(G860), .ZN(n813) );
  NAND2_X1 U890 ( .A1(n801), .A2(G55), .ZN(n802) );
  XOR2_X1 U891 ( .A(KEYINPUT81), .B(n802), .Z(n805) );
  NAND2_X1 U892 ( .A1(G67), .A2(n803), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT82), .B(n806), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G93), .A2(n807), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G80), .A2(n808), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n822) );
  XOR2_X1 U899 ( .A(n813), .B(n822), .Z(G145) );
  XOR2_X1 U900 ( .A(n822), .B(G290), .Z(n819) );
  XOR2_X1 U901 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n815) );
  XNOR2_X1 U902 ( .A(n979), .B(G288), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U904 ( .A(G166), .B(n816), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n817), .B(G305), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n819), .B(n818), .ZN(n912) );
  XNOR2_X1 U907 ( .A(n820), .B(n912), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n821), .A2(G868), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n825), .A2(n824), .ZN(G295) );
  XOR2_X1 U911 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n827) );
  NAND2_X1 U912 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XNOR2_X1 U913 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U914 ( .A1(G2090), .A2(n828), .ZN(n829) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G236), .A2(G238), .ZN(n831) );
  NAND2_X1 U919 ( .A1(G69), .A2(n831), .ZN(n832) );
  NOR2_X1 U920 ( .A1(n832), .A2(G237), .ZN(n833) );
  XNOR2_X1 U921 ( .A(n833), .B(KEYINPUT91), .ZN(n846) );
  NAND2_X1 U922 ( .A1(n846), .A2(G567), .ZN(n840) );
  NOR2_X1 U923 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U924 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U925 ( .A1(G218), .A2(n835), .ZN(n836) );
  XOR2_X1 U926 ( .A(KEYINPUT89), .B(n836), .Z(n837) );
  NAND2_X1 U927 ( .A1(G96), .A2(n837), .ZN(n838) );
  XNOR2_X1 U928 ( .A(KEYINPUT90), .B(n838), .ZN(n847) );
  NAND2_X1 U929 ( .A1(n847), .A2(G2106), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n848) );
  NAND2_X1 U931 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n848), .A2(n841), .ZN(n845) );
  NAND2_X1 U933 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U936 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n848), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U947 ( .A(n851), .B(G2100), .Z(n853) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U950 ( .A(G2096), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT109), .B(G2678), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(n857), .B(n856), .Z(G227) );
  XOR2_X1 U954 ( .A(G1986), .B(G1981), .Z(n859) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1971), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n869) );
  XOR2_X1 U957 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n861) );
  XNOR2_X1 U958 ( .A(G1996), .B(KEYINPUT111), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U960 ( .A(G1991), .B(G1976), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1961), .B(G1956), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT112), .B(G2474), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G124), .A2(n901), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U969 ( .A1(n900), .A2(G112), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G100), .A2(n524), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G136), .A2(n525), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U975 ( .A(n877), .B(G162), .ZN(n879) );
  XNOR2_X1 U976 ( .A(G164), .B(G160), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n895) );
  XNOR2_X1 U978 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G106), .A2(n524), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G142), .A2(n525), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(KEYINPUT45), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G118), .A2(n900), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G130), .A2(n901), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(KEYINPUT115), .B(n891), .Z(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n908) );
  NAND2_X1 U993 ( .A1(G103), .A2(n524), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G139), .A2(n525), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G115), .A2(n900), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G127), .A2(n901), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n964) );
  XNOR2_X1 U1001 ( .A(n964), .B(n954), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT116), .B(n912), .Z(n915) );
  XNOR2_X1 U1006 ( .A(n913), .B(G286), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1008 ( .A(n992), .B(G171), .Z(n916) );
  XNOR2_X1 U1009 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n920), .ZN(n921) );
  AND2_X1 U1014 ( .A1(G319), .A2(n921), .ZN(n923) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1019 ( .A(G1348), .B(KEYINPUT59), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(G4), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G1956), .B(G20), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G1981), .B(G6), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1025 ( .A(KEYINPUT123), .B(G1341), .Z(n929) );
  XNOR2_X1 U1026 ( .A(G19), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT60), .B(n932), .ZN(n944) );
  XOR2_X1 U1029 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n939) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(G24), .B(G1986), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1033 ( .A(G1976), .B(KEYINPUT124), .Z(n935) );
  XNOR2_X1 U1034 ( .A(G23), .B(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n939), .B(n938), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G1961), .B(KEYINPUT122), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(G5), .B(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G21), .B(G1966), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1043 ( .A(KEYINPUT61), .B(n947), .Z(n948) );
  NOR2_X1 U1044 ( .A1(G16), .A2(n948), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT126), .B(n949), .Z(n950) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n950), .ZN(n978) );
  XOR2_X1 U1047 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT51), .B(n953), .Z(n963) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G2084), .B(G160), .Z(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n971) );
  XOR2_X1 U1056 ( .A(G2072), .B(n964), .Z(n966) );
  XOR2_X1 U1057 ( .A(G164), .B(G2078), .Z(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(n967), .B(KEYINPUT50), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(n972), .B(KEYINPUT52), .ZN(n974) );
  INV_X1 U1063 ( .A(KEYINPUT55), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(G29), .A2(n975), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT117), .B(n976), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n1028) );
  XOR2_X1 U1068 ( .A(KEYINPUT56), .B(G16), .Z(n1003) );
  XNOR2_X1 U1069 ( .A(n979), .B(G1956), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n991) );
  XNOR2_X1 U1072 ( .A(n984), .B(KEYINPUT121), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(n985), .B(G1348), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G303), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n1001) );
  XNOR2_X1 U1078 ( .A(G301), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(n992), .B(G1341), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n999) );
  XOR2_X1 U1081 ( .A(G168), .B(G1966), .Z(n995) );
  NOR2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n997), .Z(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1086 ( .A1(n1003), .A2(n1002), .ZN(n1026) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1019) );
  XOR2_X1 U1088 ( .A(G1991), .B(G25), .Z(n1004) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(G28), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(KEYINPUT118), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(n1006), .B(G27), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G32), .B(G1996), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(KEYINPUT119), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G2067), .B(G26), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G33), .B(G2072), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1016), .B(KEYINPUT53), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(n1017), .B(KEYINPUT120), .ZN(n1018) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(KEYINPUT54), .B(G2084), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(G34), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT55), .B(n1023), .Z(n1024) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1029), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

