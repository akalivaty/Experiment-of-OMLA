

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597;

  XOR2_X1 U323 ( .A(KEYINPUT123), .B(n463), .Z(n590) );
  NOR2_X2 U324 ( .A1(n491), .A2(n566), .ZN(n463) );
  INV_X1 U325 ( .A(G22GAT), .ZN(n433) );
  XNOR2_X1 U326 ( .A(G155GAT), .B(KEYINPUT91), .ZN(n408) );
  XNOR2_X1 U327 ( .A(n420), .B(n291), .ZN(n421) );
  XNOR2_X1 U328 ( .A(n348), .B(n347), .ZN(n349) );
  INV_X1 U329 ( .A(G197GAT), .ZN(n347) );
  XNOR2_X1 U330 ( .A(n487), .B(KEYINPUT38), .ZN(n517) );
  NOR2_X1 U331 ( .A1(n533), .A2(n502), .ZN(n487) );
  AND2_X1 U332 ( .A1(G225GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U333 ( .A(KEYINPUT98), .B(n469), .Z(n292) );
  XNOR2_X1 U334 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n358) );
  NOR2_X1 U335 ( .A1(n475), .A2(n474), .ZN(n476) );
  INV_X1 U336 ( .A(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U337 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U338 ( .A(n410), .B(n409), .ZN(n411) );
  INV_X1 U339 ( .A(KEYINPUT48), .ZN(n403) );
  XNOR2_X1 U340 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U341 ( .A(n412), .B(n411), .ZN(n441) );
  XNOR2_X1 U342 ( .A(n403), .B(KEYINPUT64), .ZN(n404) );
  NOR2_X1 U343 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U344 ( .A(n350), .B(n349), .ZN(n355) );
  XNOR2_X1 U345 ( .A(n422), .B(n421), .ZN(n430) );
  XNOR2_X1 U346 ( .A(n485), .B(KEYINPUT41), .ZN(n577) );
  XOR2_X1 U347 ( .A(n445), .B(n444), .Z(n490) );
  INV_X1 U348 ( .A(G204GAT), .ZN(n464) );
  XNOR2_X1 U349 ( .A(KEYINPUT96), .B(n478), .ZN(n534) );
  XNOR2_X1 U350 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n488) );
  XNOR2_X1 U352 ( .A(n467), .B(n466), .ZN(G1353GAT) );
  XNOR2_X1 U353 ( .A(n489), .B(n488), .ZN(G1330GAT) );
  XOR2_X1 U354 ( .A(G176GAT), .B(G183GAT), .Z(n294) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U357 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n296) );
  XNOR2_X1 U358 ( .A(G190GAT), .B(KEYINPUT85), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U360 ( .A(n298), .B(n297), .Z(n460) );
  XOR2_X1 U361 ( .A(KEYINPUT90), .B(G218GAT), .Z(n300) );
  XNOR2_X1 U362 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U364 ( .A(G197GAT), .B(n301), .Z(n444) );
  XNOR2_X1 U365 ( .A(n460), .B(n444), .ZN(n308) );
  XNOR2_X1 U366 ( .A(G92GAT), .B(G64GAT), .ZN(n311) );
  INV_X1 U367 ( .A(n311), .ZN(n314) );
  XOR2_X1 U368 ( .A(KEYINPUT97), .B(G204GAT), .Z(n303) );
  XNOR2_X1 U369 ( .A(G36GAT), .B(G8GAT), .ZN(n302) );
  XNOR2_X1 U370 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U371 ( .A(n314), .B(n304), .Z(n306) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U373 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U374 ( .A(n308), .B(n307), .ZN(n537) );
  INV_X1 U375 ( .A(G57GAT), .ZN(n309) );
  NAND2_X1 U376 ( .A1(n309), .A2(G148GAT), .ZN(n313) );
  INV_X1 U377 ( .A(G148GAT), .ZN(n310) );
  NAND2_X1 U378 ( .A1(n310), .A2(G57GAT), .ZN(n312) );
  NAND2_X1 U379 ( .A1(n313), .A2(n312), .ZN(n413) );
  NAND2_X1 U380 ( .A1(n413), .A2(n311), .ZN(n317) );
  AND2_X1 U381 ( .A1(n313), .A2(n312), .ZN(n315) );
  NAND2_X1 U382 ( .A1(n315), .A2(n314), .ZN(n316) );
  NAND2_X1 U383 ( .A1(n317), .A2(n316), .ZN(n319) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U385 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U386 ( .A(KEYINPUT13), .B(KEYINPUT31), .Z(n321) );
  XNOR2_X1 U387 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U389 ( .A(n323), .B(n322), .ZN(n330) );
  INV_X1 U390 ( .A(n330), .ZN(n328) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G71GAT), .Z(n449) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U393 ( .A(G120GAT), .B(G176GAT), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U395 ( .A(n449), .B(n326), .Z(n329) );
  INV_X1 U396 ( .A(n329), .ZN(n327) );
  NAND2_X1 U397 ( .A1(n328), .A2(n327), .ZN(n332) );
  NAND2_X1 U398 ( .A1(n330), .A2(n329), .ZN(n331) );
  NAND2_X1 U399 ( .A1(n332), .A2(n331), .ZN(n334) );
  INV_X1 U400 ( .A(KEYINPUT72), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U402 ( .A(G78GAT), .B(G204GAT), .Z(n336) );
  XNOR2_X1 U403 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U404 ( .A(n336), .B(n335), .ZN(n436) );
  XNOR2_X1 U405 ( .A(n436), .B(KEYINPUT70), .ZN(n337) );
  XNOR2_X2 U406 ( .A(n338), .B(n337), .ZN(n485) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT7), .Z(n340) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(G36GAT), .ZN(n339) );
  XNOR2_X1 U409 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U410 ( .A(KEYINPUT8), .B(n341), .Z(n384) );
  XOR2_X1 U411 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G113GAT), .ZN(n342) );
  XNOR2_X1 U413 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n384), .B(n344), .ZN(n357) );
  XOR2_X1 U415 ( .A(G1GAT), .B(G8GAT), .Z(n346) );
  XNOR2_X1 U416 ( .A(G22GAT), .B(G15GAT), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n360) );
  XNOR2_X1 U418 ( .A(G141GAT), .B(n360), .ZN(n350) );
  XOR2_X1 U419 ( .A(G29GAT), .B(G43GAT), .Z(n348) );
  XOR2_X1 U420 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n352) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U422 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U423 ( .A(KEYINPUT66), .B(n353), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n583) );
  NAND2_X1 U426 ( .A1(n577), .A2(n583), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n379) );
  XOR2_X1 U428 ( .A(n360), .B(KEYINPUT79), .Z(n362) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U431 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n364) );
  XNOR2_X1 U432 ( .A(KEYINPUT13), .B(KEYINPUT78), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n376) );
  XOR2_X1 U434 ( .A(G78GAT), .B(G155GAT), .Z(n366) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n368) );
  XNOR2_X1 U438 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U440 ( .A(G57GAT), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U441 ( .A(G183GAT), .B(G71GAT), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U443 ( .A(n372), .B(n371), .Z(n373) );
  XNOR2_X1 U444 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U445 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n557) );
  NAND2_X1 U447 ( .A1(n379), .A2(n557), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n380), .B(KEYINPUT115), .ZN(n395) );
  XOR2_X1 U449 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n382) );
  XNOR2_X1 U450 ( .A(G99GAT), .B(KEYINPUT10), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT9), .B(G92GAT), .Z(n386) );
  XNOR2_X1 U454 ( .A(G162GAT), .B(G106GAT), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U456 ( .A(G29GAT), .B(G85GAT), .Z(n414) );
  XOR2_X1 U457 ( .A(n414), .B(G218GAT), .Z(n388) );
  XOR2_X1 U458 ( .A(G43GAT), .B(G134GAT), .Z(n456) );
  XNOR2_X1 U459 ( .A(G190GAT), .B(n456), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U461 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U462 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U463 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n494) );
  NAND2_X1 U465 ( .A1(n395), .A2(n494), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n396), .B(KEYINPUT47), .ZN(n402) );
  XOR2_X1 U467 ( .A(KEYINPUT36), .B(KEYINPUT105), .Z(n397) );
  XNOR2_X1 U468 ( .A(n494), .B(n397), .ZN(n594) );
  NOR2_X1 U469 ( .A1(n557), .A2(n594), .ZN(n398) );
  XNOR2_X1 U470 ( .A(KEYINPUT45), .B(n398), .ZN(n399) );
  NAND2_X1 U471 ( .A1(n399), .A2(n485), .ZN(n400) );
  NOR2_X1 U472 ( .A1(n400), .A2(n583), .ZN(n401) );
  NOR2_X1 U473 ( .A1(n402), .A2(n401), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n547) );
  NAND2_X1 U475 ( .A1(n537), .A2(n547), .ZN(n407) );
  XOR2_X1 U476 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n406) );
  XNOR2_X1 U477 ( .A(n407), .B(n406), .ZN(n431) );
  XNOR2_X1 U478 ( .A(n408), .B(KEYINPUT2), .ZN(n412) );
  XNOR2_X1 U479 ( .A(G141GAT), .B(G162GAT), .ZN(n410) );
  XOR2_X1 U480 ( .A(n414), .B(n413), .Z(n416) );
  XNOR2_X1 U481 ( .A(G1GAT), .B(G134GAT), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U483 ( .A(n441), .B(n417), .Z(n422) );
  XOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n419) );
  XNOR2_X1 U485 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U487 ( .A(KEYINPUT0), .B(G127GAT), .Z(n424) );
  XNOR2_X1 U488 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U490 ( .A(G113GAT), .B(n425), .Z(n457) );
  XOR2_X1 U491 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U492 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n457), .B(n428), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n478) );
  NOR2_X1 U496 ( .A1(n431), .A2(n534), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n432), .B(KEYINPUT65), .ZN(n491) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XOR2_X1 U499 ( .A(G148GAT), .B(KEYINPUT24), .Z(n438) );
  XNOR2_X1 U500 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U502 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U503 ( .A(G50GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT82), .B(KEYINPUT86), .Z(n447) );
  XNOR2_X1 U506 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U508 ( .A(n448), .B(KEYINPUT83), .Z(n451) );
  XNOR2_X1 U509 ( .A(G15GAT), .B(n449), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT84), .B(KEYINPUT87), .Z(n453) );
  NAND2_X1 U512 ( .A1(G227GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U514 ( .A(n455), .B(n454), .Z(n459) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(n539) );
  INV_X1 U518 ( .A(n539), .ZN(n549) );
  NAND2_X1 U519 ( .A1(n490), .A2(n549), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT26), .ZN(n566) );
  INV_X1 U521 ( .A(n590), .ZN(n595) );
  OR2_X1 U522 ( .A1(n595), .A2(n485), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n465) );
  XOR2_X1 U524 ( .A(n537), .B(KEYINPUT27), .Z(n473) );
  INV_X1 U525 ( .A(n473), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n534), .A2(n468), .ZN(n546) );
  XNOR2_X1 U527 ( .A(n490), .B(KEYINPUT28), .ZN(n552) );
  NOR2_X1 U528 ( .A1(n546), .A2(n552), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n549), .B(KEYINPUT89), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n292), .A2(n470), .ZN(n480) );
  AND2_X1 U531 ( .A1(n539), .A2(n537), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n490), .A2(n471), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n472), .Z(n475) );
  NOR2_X1 U534 ( .A1(n566), .A2(n473), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT99), .B(n476), .Z(n477) );
  NOR2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n479) );
  XOR2_X1 U537 ( .A(n481), .B(KEYINPUT100), .Z(n500) );
  AND2_X1 U538 ( .A1(n557), .A2(n500), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT106), .B(n482), .Z(n483) );
  NOR2_X1 U540 ( .A1(n594), .A2(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n484), .ZN(n533) );
  NAND2_X1 U542 ( .A1(n485), .A2(n583), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT74), .ZN(n502) );
  NAND2_X1 U544 ( .A1(n539), .A2(n517), .ZN(n489) );
  NOR2_X1 U545 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U546 ( .A(n492), .B(KEYINPUT55), .ZN(n493) );
  NOR2_X2 U547 ( .A1(n549), .A2(n493), .ZN(n581) );
  INV_X1 U548 ( .A(n494), .ZN(n574) );
  NAND2_X1 U549 ( .A1(n581), .A2(n574), .ZN(n498) );
  XOR2_X1 U550 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n496) );
  INV_X1 U551 ( .A(G190GAT), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U553 ( .A(n498), .B(n497), .ZN(G1351GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n505) );
  NOR2_X1 U555 ( .A1(n557), .A2(n574), .ZN(n499) );
  XNOR2_X1 U556 ( .A(KEYINPUT16), .B(n499), .ZN(n501) );
  NAND2_X1 U557 ( .A1(n501), .A2(n500), .ZN(n520) );
  NOR2_X1 U558 ( .A1(n502), .A2(n520), .ZN(n503) );
  XOR2_X1 U559 ( .A(KEYINPUT101), .B(n503), .Z(n510) );
  NAND2_X1 U560 ( .A1(n510), .A2(n534), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U562 ( .A(G1GAT), .B(n506), .Z(G1324GAT) );
  NAND2_X1 U563 ( .A1(n510), .A2(n537), .ZN(n507) );
  XNOR2_X1 U564 ( .A(n507), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .Z(n509) );
  NAND2_X1 U566 ( .A1(n510), .A2(n539), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n512) );
  NAND2_X1 U569 ( .A1(n510), .A2(n552), .ZN(n511) );
  XNOR2_X1 U570 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(n513), .ZN(G1327GAT) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n515) );
  NAND2_X1 U573 ( .A1(n517), .A2(n534), .ZN(n514) );
  XNOR2_X1 U574 ( .A(n515), .B(n514), .ZN(G1328GAT) );
  NAND2_X1 U575 ( .A1(n517), .A2(n537), .ZN(n516) );
  XNOR2_X1 U576 ( .A(n516), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n517), .A2(n552), .ZN(n518) );
  XNOR2_X1 U578 ( .A(n518), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n522) );
  INV_X1 U580 ( .A(n583), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n519), .A2(n577), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n532), .A2(n520), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n529), .A2(n534), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U585 ( .A(n523), .B(KEYINPUT42), .Z(n525) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(G1332GAT) );
  NAND2_X1 U588 ( .A1(n529), .A2(n537), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n539), .A2(n529), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n531) );
  NAND2_X1 U594 ( .A1(n529), .A2(n552), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1335GAT) );
  XOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT111), .Z(n536) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n534), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n541), .A2(n537), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n539), .A2(n541), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n541), .A2(n552), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1339GAT) );
  INV_X1 U609 ( .A(n546), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n565) );
  NOR2_X1 U611 ( .A1(n549), .A2(n565), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(n550), .Z(n551) );
  NOR2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n561), .A2(n583), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n555) );
  NAND2_X1 U617 ( .A1(n561), .A2(n577), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U619 ( .A(G120GAT), .B(n556), .Z(G1341GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n559) );
  INV_X1 U621 ( .A(n557), .ZN(n589) );
  NAND2_X1 U622 ( .A1(n561), .A2(n589), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U624 ( .A(G127GAT), .B(n560), .Z(G1342GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n563) );
  NAND2_X1 U626 ( .A1(n561), .A2(n574), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(G134GAT), .B(n564), .Z(G1343GAT) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n583), .A2(n573), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G141GAT), .B(n567), .ZN(G1344GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n569) );
  NAND2_X1 U633 ( .A1(n573), .A2(n577), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G148GAT), .B(n570), .ZN(G1345GAT) );
  NAND2_X1 U636 ( .A1(n589), .A2(n573), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT120), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G155GAT), .B(n572), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U641 ( .A1(n583), .A2(n581), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G169GAT), .B(n576), .ZN(G1348GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n579) );
  NAND2_X1 U644 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(G176GAT), .B(n580), .ZN(G1349GAT) );
  NAND2_X1 U647 ( .A1(n589), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U649 ( .A1(n590), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT124), .ZN(n586) );
  INV_X1 U651 ( .A(KEYINPUT60), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(G211GAT), .B(n593), .ZN(G1354GAT) );
  NOR2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U660 ( .A(KEYINPUT62), .B(n596), .Z(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

