//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n455), .A2(KEYINPUT67), .A3(G567), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n466), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n465), .A2(KEYINPUT68), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n470), .B1(new_n479), .B2(G2105), .ZN(G160));
  NOR2_X1   g055(.A1(new_n474), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n466), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT69), .B1(new_n474), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n465), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n466), .C1(new_n472), .C2(new_n473), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n491), .A2(new_n495), .B1(KEYINPUT4), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n505), .B2(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT71), .B(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n511), .B2(new_n513), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n506), .A2(new_n516), .A3(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n522));
  AND3_X1   g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n514), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n514), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT73), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(KEYINPUT73), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n505), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n518), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n514), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n518), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n509), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n514), .A2(G91), .B1(new_n559), .B2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G299));
  OR2_X1    g136(.A1(new_n503), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(G87), .A2(new_n514), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n518), .A2(G49), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n564), .A2(KEYINPUT75), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(KEYINPUT75), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(G288));
  AND3_X1   g142(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT6), .B1(new_n512), .B2(G651), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n503), .B(G86), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(G48), .B(G543), .C1(new_n568), .C2(new_n569), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OR2_X1    g151(.A1(KEYINPUT5), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(KEYINPUT5), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n572), .A2(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n514), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n505), .C2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(new_n514), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n505), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI21_X1  g170(.A(G543), .B1(new_n568), .B2(new_n569), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g177(.A(new_n601), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n556), .A2(new_n560), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(G860), .B2(new_n609), .ZN(G148));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n547), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n614), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n481), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n483), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n466), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT81), .B(G2096), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n465), .A2(new_n468), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(KEYINPUT80), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(KEYINPUT80), .B2(new_n628), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n623), .B(new_n630), .C1(new_n631), .C2(new_n629), .ZN(G156));
  INV_X1    g207(.A(G14), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(G2438), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n634), .A2(KEYINPUT83), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n634), .A2(KEYINPUT83), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(new_n636), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n643), .A3(new_n641), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n646), .B2(KEYINPUT14), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT85), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G1341), .ZN(new_n659));
  INV_X1    g234(.A(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n633), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n655), .A3(new_n661), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n666), .C2(new_n667), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n666), .A2(new_n667), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n669), .A2(new_n676), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(new_n668), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n672), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G1986), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1961), .B(G1966), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n692), .B2(new_n696), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n690), .B(KEYINPUT19), .ZN(new_n701));
  INV_X1    g276(.A(new_n696), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n694), .A2(new_n695), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n689), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n699), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(new_n697), .ZN(new_n709));
  INV_X1    g284(.A(new_n706), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT89), .ZN(new_n711));
  INV_X1    g286(.A(G1981), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n712), .B1(new_n707), .B2(new_n711), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n688), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(new_n711), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G1981), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n721), .A2(G1986), .A3(new_n713), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n716), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n687), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n714), .A2(new_n715), .A3(new_n688), .ZN(new_n726));
  AOI21_X1  g301(.A(G1986), .B1(new_n721), .B2(new_n713), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(new_n686), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(new_n730), .ZN(G229));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G6), .ZN(new_n733));
  INV_X1    g308(.A(G305), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT32), .B(G1981), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n732), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n732), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1971), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n732), .A2(G23), .ZN(new_n742));
  INV_X1    g317(.A(G288), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n732), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT33), .B(G1976), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n738), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT34), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n481), .A2(G131), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n483), .A2(G119), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n466), .A2(G107), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G25), .B(new_n755), .S(G29), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT35), .B(G1991), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n732), .A2(G24), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G290), .B2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n758), .B1(new_n760), .B2(new_n688), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n688), .B2(new_n760), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n763), .B(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G105), .B2(new_n468), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n771));
  AOI22_X1  g346(.A1(G129), .A2(new_n483), .B1(new_n481), .B2(G141), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G29), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT27), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1996), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(G1996), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n608), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT93), .B(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n781), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n732), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n732), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT98), .Z(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(G1961), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n732), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n777), .A2(G33), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n481), .A2(G139), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT25), .Z(new_n801));
  AOI22_X1  g376(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n466), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n804), .B2(new_n777), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G19), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n548), .B2(G16), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n805), .A2(G2072), .B1(G1341), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(G2072), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n732), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n732), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(G1966), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n792), .A2(new_n796), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n777), .A2(G35), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G162), .B2(new_n777), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT29), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT24), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n777), .B1(new_n817), .B2(G34), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(G34), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G160), .B2(G29), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n816), .A2(G2090), .B1(G2084), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G2084), .B2(new_n820), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT30), .B(G28), .ZN(new_n823));
  OR2_X1    g398(.A1(KEYINPUT31), .A2(G11), .ZN(new_n824));
  NAND2_X1  g399(.A1(KEYINPUT31), .A2(G11), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n823), .A2(new_n777), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n826), .B1(new_n777), .B2(new_n621), .C1(new_n807), .C2(G1341), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n811), .A2(G1966), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n777), .A2(G26), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT94), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT28), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n481), .A2(G140), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n483), .A2(G128), .ZN(new_n833));
  OR2_X1    g408(.A1(G104), .A2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n831), .B1(new_n837), .B2(new_n777), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G2067), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n827), .A2(new_n828), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n777), .A2(G27), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G164), .B2(new_n777), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G2078), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n816), .B2(G2090), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n822), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NOR4_X1   g420(.A1(new_n787), .A2(new_n791), .A3(new_n813), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n766), .A2(new_n846), .ZN(G150));
  INV_X1    g422(.A(G150), .ZN(G311));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n509), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n505), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n514), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n854), .A2(new_n860), .A3(new_n855), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n854), .B2(new_n855), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n547), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n854), .A2(new_n860), .A3(new_n855), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n548), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n608), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n870));
  XOR2_X1   g445(.A(new_n869), .B(new_n870), .Z(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n859), .B1(new_n873), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(KEYINPUT106), .B(G37), .ZN(new_n877));
  INV_X1    g452(.A(new_n775), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n837), .B1(new_n878), .B2(new_n773), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n774), .A2(new_n775), .A3(new_n836), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n481), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n483), .A2(G130), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(KEYINPUT105), .B1(new_n884), .B2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(KEYINPUT105), .B2(new_n883), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n879), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n879), .B2(new_n880), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n490), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n492), .B1(new_n465), .B2(new_n494), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n501), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n804), .B(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n755), .B(new_n625), .Z(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n891), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G160), .B(new_n621), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n487), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n889), .A2(new_n906), .A3(new_n890), .A4(new_n907), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n877), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g491(.A1(G290), .A2(new_n734), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n586), .A2(G305), .A3(new_n587), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G288), .B(G303), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n614), .A2(new_n867), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n613), .A2(new_n866), .A3(new_n863), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n600), .A2(G299), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n605), .A2(new_n591), .A3(new_n599), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n925), .A3(new_n926), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n932), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n932), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n924), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g518(.A(new_n924), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n932), .A2(new_n937), .A3(new_n938), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n946), .A3(G868), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n856), .B2(new_n611), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n941), .A2(new_n946), .A3(KEYINPUT107), .A4(G868), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G295));
  AND2_X1   g529(.A1(new_n949), .A2(new_n951), .ZN(G331));
  AOI21_X1  g530(.A(new_n934), .B1(new_n928), .B2(new_n929), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n935), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n931), .A2(KEYINPUT110), .A3(new_n934), .ZN(new_n959));
  OAI21_X1  g534(.A(G286), .B1(new_n539), .B2(new_n540), .ZN(new_n960));
  INV_X1    g535(.A(new_n540), .ZN(new_n961));
  NAND3_X1  g536(.A1(G168), .A2(new_n961), .A3(new_n538), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n863), .A2(new_n866), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n867), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n958), .A2(new_n959), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n931), .A3(new_n963), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n944), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n936), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n924), .A3(new_n967), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n877), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g549(.A(G37), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n924), .B1(new_n971), .B2(new_n967), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n974), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n969), .A2(new_n981), .A3(new_n877), .A4(new_n972), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n903), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n989), .B(new_n470), .C1(new_n479), .C2(G2105), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n836), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n776), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n991), .A2(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n776), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n992), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n755), .B(new_n757), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n991), .ZN(new_n1006));
  XNOR2_X1  g581(.A(G290), .B(G1986), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n903), .A2(new_n987), .A3(new_n990), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n563), .B(G1976), .C1(new_n565), .C2(new_n566), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(G8), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n570), .A2(new_n571), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n573), .B(KEYINPUT76), .ZN(new_n1014));
  OAI21_X1  g589(.A(G61), .B1(new_n507), .B2(new_n508), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n505), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n580), .A2(new_n712), .A3(new_n571), .A4(new_n570), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1023), .A2(G8), .A3(new_n1009), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1009), .A2(new_n1029), .A3(G8), .A4(new_n1010), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1012), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1012), .A2(new_n1027), .A3(new_n1033), .A4(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT55), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n479), .A2(G2105), .ZN(new_n1039));
  INV_X1    g614(.A(new_n470), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G40), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n501), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n895), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT113), .B1(new_n1043), .B2(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n987), .B1(new_n497), .B2(new_n501), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1041), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1971), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1041), .B1(new_n1045), .B2(KEYINPUT50), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n903), .A2(new_n1053), .A3(new_n987), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G2090), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(new_n1038), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1050), .A3(new_n990), .ZN(new_n1059));
  INV_X1    g634(.A(G1971), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1053), .B(new_n987), .C1(new_n497), .C2(new_n501), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n990), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n903), .A2(new_n987), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g639(.A(G2090), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1059), .A2(new_n1060), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1037), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G168), .A2(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(new_n1047), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n990), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2084), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1052), .A2(new_n1054), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1069), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1035), .A2(new_n1057), .A3(new_n1068), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1068), .A2(new_n1057), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1035), .A4(new_n1078), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1037), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1031), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1078), .A3(new_n1089), .A4(new_n1057), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1009), .A2(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n743), .A2(new_n1028), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1027), .A2(new_n1096), .B1(new_n712), .B2(new_n734), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1057), .A2(new_n1031), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G2078), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1058), .A2(new_n1099), .A3(new_n1050), .A4(new_n990), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1055), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n988), .A2(new_n1041), .A3(new_n1071), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1035), .A2(new_n1107), .A3(new_n1057), .A4(new_n1068), .ZN(new_n1108));
  OAI211_X1 g683(.A(G168), .B(new_n1077), .C1(new_n1104), .C2(G1966), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(G168), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1108), .B1(new_n1115), .B2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1098), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1093), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n605), .B(KEYINPUT57), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1049), .A2(new_n1050), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1053), .B1(new_n903), .B2(new_n987), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(new_n1062), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1121), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1123), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1009), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n903), .A2(KEYINPUT119), .A3(new_n990), .A4(new_n987), .ZN(new_n1132));
  AOI21_X1  g707(.A(G2067), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1348), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n608), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT120), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1128), .B(new_n1138), .C1(new_n1129), .C2(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1129), .B2(new_n1127), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n608), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n600), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1147), .B2(new_n1135), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1129), .A2(new_n1127), .A3(new_n1141), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  NAND3_X1  g726(.A1(new_n1131), .A2(new_n1132), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1049), .A2(new_n995), .A3(new_n1050), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n548), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n1155), .B2(KEYINPUT59), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n547), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT121), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT59), .B1(new_n1157), .B2(KEYINPUT121), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1157), .A2(KEYINPUT121), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n1158), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1140), .B1(new_n1150), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(G301), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1070), .A2(KEYINPUT123), .A3(new_n990), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n988), .B2(new_n1041), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1170), .A2(new_n1172), .A3(new_n1050), .A4(new_n1105), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1103), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1174), .B2(G171), .ZN(new_n1175));
  AOI211_X1 g750(.A(KEYINPUT124), .B(G301), .C1(new_n1103), .C2(new_n1173), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1174), .A2(G171), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1166), .B1(new_n1178), .B2(new_n1107), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1035), .A2(new_n1057), .A3(new_n1068), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1115), .A4(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1008), .B1(new_n1120), .B2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n998), .A2(KEYINPUT46), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n776), .A2(new_n994), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n992), .A2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1188), .B(new_n1190), .C1(KEYINPUT46), .C2(new_n998), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1191), .A2(KEYINPUT47), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(KEYINPUT47), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1005), .A2(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n757), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n755), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1002), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n837), .A2(new_n993), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1003), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1183), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g776(.A1(G227), .A2(new_n463), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n663), .B2(new_n664), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n725), .A2(new_n730), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n725), .A2(new_n1204), .A3(new_n730), .A4(KEYINPUT126), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n983), .A2(new_n1207), .A3(new_n915), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1209), .A2(KEYINPUT127), .ZN(new_n1210));
  AND2_X1   g784(.A1(new_n915), .A2(new_n1208), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1212));
  NAND4_X1  g786(.A1(new_n1211), .A2(new_n1212), .A3(new_n983), .A4(new_n1207), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n1210), .A2(new_n1213), .ZN(G308));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(G225));
endmodule


