//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT83), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n191), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n189), .B2(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G104), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G104), .A3(new_n210), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n211), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n210), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n195), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G128), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n191), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n190), .A2(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n231), .B1(new_n203), .B2(new_n207), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n238), .B2(G134), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n236), .B2(G137), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT11), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT67), .B(G131), .C1(new_n241), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(KEYINPUT11), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n240), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT66), .B(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n237), .A4(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n247), .A3(new_n237), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT67), .B1(new_n251), .B2(G131), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n235), .A2(KEYINPUT12), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT85), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n235), .A2(new_n257), .A3(KEYINPUT12), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n235), .A2(new_n254), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n225), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n266), .A2(new_n218), .B1(G104), .B2(new_n210), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n219), .A2(new_n217), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n265), .B(G101), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n203), .A2(new_n270), .B1(new_n231), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G101), .B1(new_n267), .B2(new_n268), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n228), .A2(G128), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT68), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n231), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n208), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n274), .A2(new_n276), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n245), .A2(new_n249), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n252), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n264), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT84), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT84), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n264), .A2(new_n282), .A3(new_n287), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G110), .B(G140), .ZN(new_n290));
  INV_X1    g104(.A(G953), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n291), .A2(G227), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n290), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n262), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n219), .A2(new_n217), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n215), .B1(new_n297), .B2(new_n214), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n269), .A2(new_n273), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n301));
  OAI22_X1  g115(.A1(new_n299), .A2(new_n300), .B1(new_n232), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT10), .B1(new_n209), .B2(new_n224), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n254), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n294), .B1(new_n289), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n187), .B(new_n188), .C1(new_n295), .C2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n293), .B1(new_n286), .B2(new_n288), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n304), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n262), .A2(new_n289), .ZN(new_n309));
  OAI211_X1 g123(.A(G469), .B(new_n308), .C1(new_n309), .C2(new_n294), .ZN(new_n310));
  NAND2_X1  g124(.A1(G469), .A2(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G214), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n318));
  INV_X1    g132(.A(G113), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT70), .B1(KEYINPUT2), .B2(G113), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT2), .A2(G113), .ZN(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G119), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n322), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n321), .ZN(new_n328));
  NOR3_X1   g142(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT71), .A3(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n327), .A2(new_n276), .A3(new_n334), .A4(new_n269), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(G116), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT86), .A4(G116), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n336), .A2(G113), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n224), .A2(new_n333), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n327), .A2(new_n334), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n269), .B1(new_n296), .B2(new_n298), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n347), .B(new_n344), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT6), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n347), .B1(new_n335), .B2(new_n344), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n315), .B(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n354), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n352), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n273), .A2(G125), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n232), .B2(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n291), .A2(G224), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT88), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT89), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n360), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n347), .B(KEYINPUT8), .ZN(new_n368));
  AND4_X1   g182(.A1(new_n333), .A2(new_n343), .A3(new_n223), .A4(new_n220), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n343), .A2(new_n333), .B1(new_n223), .B2(new_n220), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n359), .B(new_n372), .C1(new_n232), .C2(G125), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n374), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n352), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n371), .A2(new_n374), .A3(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n366), .A2(new_n367), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n367), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n364), .B1(new_n355), .B2(new_n357), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n188), .B1(new_n386), .B2(new_n378), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n314), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G221), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n392), .B2(new_n188), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n312), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G472), .A2(G902), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT31), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n350), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n273), .B1(new_n283), .B2(new_n252), .ZN(new_n400));
  INV_X1    g214(.A(new_n237), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n236), .A2(G137), .ZN(new_n402));
  OAI21_X1  g216(.A(G131), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n249), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n281), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n327), .A2(new_n334), .A3(KEYINPUT73), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n399), .A2(new_n400), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT74), .B(KEYINPUT27), .Z(new_n410));
  NOR2_X1   g224(.A1(G237), .A2(G953), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G210), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT26), .B(G101), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT69), .B1(new_n232), .B2(new_n404), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n281), .A2(new_n419), .A3(new_n249), .A4(new_n403), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n400), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n405), .B2(new_n281), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n350), .B1(new_n424), .B2(new_n400), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n423), .A2(KEYINPUT72), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT72), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n397), .B(new_n417), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n408), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n350), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n421), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n433), .B2(new_n408), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n416), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n425), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n423), .A2(KEYINPUT72), .A3(new_n425), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n397), .B1(new_n441), .B2(new_n417), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n396), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT32), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n417), .B1(new_n426), .B2(new_n427), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT31), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n435), .A3(new_n428), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n444), .A2(G472), .A3(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n399), .A2(new_n407), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n400), .A2(new_n406), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT75), .A3(new_n408), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(KEYINPUT28), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n458), .B(new_n416), .C1(new_n429), .C2(new_n408), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n415), .B1(new_n441), .B2(new_n408), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n399), .A2(new_n407), .ZN(new_n462));
  INV_X1    g276(.A(new_n452), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n421), .B2(new_n432), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n415), .B(new_n430), .C1(new_n464), .C2(new_n429), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n460), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G472), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n445), .A2(new_n450), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G217), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(G234), .B2(new_n188), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n204), .B2(G119), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n338), .A2(KEYINPUT76), .A3(G128), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n476), .A2(new_n477), .B1(G119), .B2(new_n204), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT24), .B(G110), .Z(new_n479));
  OR3_X1    g293(.A1(new_n478), .A2(KEYINPUT80), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT80), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT77), .B1(new_n338), .B2(G128), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n482), .A2(KEYINPUT23), .B1(new_n338), .B2(G128), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(KEYINPUT23), .B2(new_n482), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n480), .B(new_n481), .C1(G110), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G125), .B(G140), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT16), .ZN(new_n487));
  INV_X1    g301(.A(G125), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n488), .A2(KEYINPUT16), .A3(G140), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(G146), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n189), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n484), .A2(G110), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n189), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n490), .A3(KEYINPUT79), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n478), .A2(new_n479), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT79), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n499), .A3(new_n189), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n492), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT22), .B(G137), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n291), .A2(G221), .A3(G234), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n503), .B(new_n504), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n492), .B(new_n505), .C1(new_n494), .C2(new_n501), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n188), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n474), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n510), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n507), .A2(new_n188), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n472), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n508), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n515), .A2(G902), .A3(new_n471), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G113), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n216), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n411), .A2(G143), .A3(G214), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(G143), .B1(new_n411), .B2(G214), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n486), .B(new_n189), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n497), .A2(new_n500), .ZN(new_n529));
  INV_X1    g343(.A(new_n248), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT17), .B(new_n530), .C1(new_n521), .C2(new_n522), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n521), .B2(new_n522), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n291), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n191), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n248), .A3(new_n520), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(KEYINPUT91), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n523), .A2(new_n538), .A3(new_n248), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT17), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n529), .B(new_n531), .C1(new_n540), .C2(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(KEYINPUT94), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n519), .B(new_n528), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n519), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n537), .A2(new_n546), .A3(new_n539), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n537), .B2(new_n539), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n486), .B1(KEYINPUT93), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n486), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n490), .B1(new_n552), .B2(G146), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n528), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT20), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT20), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n540), .A2(KEYINPUT94), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n564), .A2(new_n529), .A3(new_n542), .A4(new_n531), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n519), .B1(new_n565), .B2(new_n528), .ZN(new_n566));
  INV_X1    g380(.A(new_n544), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n188), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G475), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n571));
  INV_X1    g385(.A(G122), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(G116), .ZN(new_n573));
  INV_X1    g387(.A(G116), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(KEYINPUT95), .A3(G122), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(G116), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(KEYINPUT96), .A3(new_n577), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n210), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n576), .A2(KEYINPUT14), .B1(G116), .B2(new_n572), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(KEYINPUT14), .B2(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G107), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT97), .B1(new_n204), .B2(G143), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n191), .A3(G128), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n587), .A2(new_n589), .B1(new_n204), .B2(G143), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n236), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n583), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n582), .B(G107), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n204), .A2(G143), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(G134), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n590), .A2(new_n595), .A3(G134), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n592), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n391), .A2(new_n470), .A3(G953), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n592), .B(new_n601), .C1(new_n593), .C2(new_n599), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n602), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n188), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G952), .ZN(new_n612));
  AOI211_X1 g426(.A(G953), .B(new_n612), .C1(G234), .C2(G237), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT21), .B(G898), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT99), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n188), .B(new_n291), .C1(G234), .C2(G237), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n570), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n395), .A2(new_n469), .A3(new_n517), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AND3_X1   g434(.A1(new_n312), .A2(new_n394), .A3(new_n517), .ZN(new_n621));
  NAND2_X1  g435(.A1(KEYINPUT100), .A2(G472), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n188), .B(new_n622), .C1(new_n436), .C2(new_n442), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n448), .B2(new_n188), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n606), .A2(new_n628), .A3(new_n607), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n603), .A2(KEYINPUT33), .A3(new_n605), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n609), .A2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n608), .A2(new_n609), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n570), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n617), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n389), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  AOI22_X1  g456(.A1(new_n560), .A2(new_n562), .B1(new_n568), .B2(G475), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n617), .B(KEYINPUT101), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n367), .B1(new_n366), .B2(new_n382), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n385), .A2(new_n387), .A3(new_n384), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n313), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NAND2_X1  g466(.A1(new_n509), .A2(new_n510), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n513), .A3(new_n473), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n471), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n502), .A2(KEYINPUT102), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n502), .A2(KEYINPUT102), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n657), .B1(new_n656), .B2(new_n658), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n188), .B(new_n472), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n610), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n608), .B(new_n663), .ZN(new_n664));
  AND4_X1   g478(.A1(new_n637), .A2(new_n662), .A3(new_n664), .A4(new_n643), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n395), .A3(new_n626), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AND2_X1   g482(.A1(new_n395), .A2(new_n469), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n669), .A2(new_n662), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n616), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n613), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n644), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  NOR2_X1   g492(.A1(new_n646), .A2(new_n647), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n570), .A2(new_n611), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n680), .A2(new_n314), .A3(new_n662), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n312), .A2(new_n394), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n674), .B(KEYINPUT39), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n454), .A2(new_n456), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n188), .B1(new_n688), .B2(new_n415), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n416), .B1(new_n441), .B2(new_n408), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n445), .A2(new_n450), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n682), .A2(new_n686), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT103), .B(G143), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G45));
  INV_X1    g509(.A(new_n634), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n643), .A3(new_n675), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n670), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(new_n517), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n467), .A2(G472), .B1(new_n448), .B2(new_n449), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(new_n445), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n302), .A2(new_n303), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n287), .B1(new_n703), .B2(new_n284), .ZN(new_n704));
  INV_X1    g518(.A(new_n288), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n304), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n706), .A2(new_n293), .B1(new_n307), .B2(new_n262), .ZN(new_n707));
  OAI21_X1  g521(.A(G469), .B1(new_n707), .B2(G902), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n394), .A3(new_n306), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(KEYINPUT104), .A3(new_n306), .A4(new_n394), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n639), .A2(new_n702), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n469), .A2(new_n517), .A3(new_n711), .A4(new_n712), .ZN(new_n717));
  INV_X1    g531(.A(new_n649), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT105), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n713), .A2(new_n720), .A3(new_n649), .A4(new_n702), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND3_X1  g537(.A1(new_n711), .A2(new_n389), .A3(new_n712), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n711), .A2(new_n726), .A3(new_n389), .A4(new_n712), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n665), .A2(new_n469), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n457), .A2(new_n430), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n732), .B(new_n447), .C1(new_n733), .C2(new_n415), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n415), .B1(new_n457), .B2(new_n430), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n442), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n736), .A3(new_n428), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n396), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n448), .A2(new_n188), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G472), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n738), .A2(new_n517), .A3(new_n740), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n389), .A2(new_n570), .A3(new_n611), .A4(new_n645), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n713), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT108), .B(G122), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G24));
  NAND4_X1  g559(.A1(new_n738), .A2(new_n697), .A3(new_n662), .A4(new_n740), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n728), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT109), .B(G125), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G27));
  AND3_X1   g564(.A1(new_n383), .A2(new_n313), .A3(new_n388), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n312), .A3(new_n394), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n469), .A3(new_n517), .A4(new_n697), .ZN(new_n753));
  NOR2_X1   g567(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n754), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n702), .A2(new_n697), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT111), .B1(new_n755), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT112), .B(G131), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G33));
  NAND3_X1  g576(.A1(new_n702), .A2(new_n676), .A3(new_n752), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NOR2_X1   g578(.A1(new_n696), .A2(new_n570), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT113), .B(KEYINPUT43), .Z(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n696), .A2(new_n570), .B1(KEYINPUT113), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(new_n662), .C1(new_n624), .C2(new_n625), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n751), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n308), .B1(new_n309), .B2(new_n294), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n311), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n311), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n306), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n394), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n684), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n773), .A2(new_n791), .A3(new_n775), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n777), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND3_X1  g608(.A1(new_n697), .A2(new_n700), .A3(new_n751), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n469), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n394), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(new_n763), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n570), .A2(new_n611), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n469), .A2(new_n802), .A3(new_n662), .A4(new_n674), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n746), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n752), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n758), .B2(new_n759), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n648), .B1(new_n635), .B2(new_n644), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n626), .A3(new_n621), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n717), .B2(new_n638), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n619), .A2(new_n666), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n722), .A3(new_n730), .A4(new_n743), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n669), .B(new_n662), .C1(new_n676), .C2(new_n697), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n681), .A2(new_n314), .A3(new_n679), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n674), .B(KEYINPUT116), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n662), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n692), .A3(new_n683), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n748), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n748), .A2(new_n818), .A3(KEYINPUT52), .A4(new_n814), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n813), .A2(KEYINPUT115), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n806), .B2(new_n812), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n804), .A2(new_n752), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n763), .ZN(new_n828));
  INV_X1    g642(.A(new_n759), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n757), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n722), .A2(new_n730), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n619), .A2(new_n666), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n743), .A3(new_n714), .A4(new_n808), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n821), .A2(new_n822), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n825), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n823), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n825), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(KEYINPUT54), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n839), .B1(new_n755), .B2(new_n757), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n805), .A2(new_n845), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n846), .B(new_n812), .C1(new_n821), .C2(new_n822), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n844), .B1(KEYINPUT54), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n708), .A2(new_n306), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(new_n393), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n797), .A2(new_n798), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n673), .B1(new_n767), .B2(new_n769), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n741), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n774), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT118), .Z(new_n859));
  OR2_X1    g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n713), .A2(new_n751), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n861), .A2(new_n700), .A3(new_n673), .A4(new_n692), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n643), .A3(new_n696), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n738), .A2(new_n662), .A3(new_n740), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n713), .A3(new_n751), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n713), .A2(new_n314), .A3(new_n680), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n868), .A2(KEYINPUT120), .A3(KEYINPUT50), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(KEYINPUT120), .B2(KEYINPUT50), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT51), .B1(new_n860), .B2(new_n871), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n612), .B(G953), .C1(new_n862), .C2(new_n636), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT48), .ZN(new_n874));
  INV_X1    g688(.A(new_n702), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT121), .B(new_n874), .C1(new_n865), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n728), .A2(new_n741), .A3(new_n856), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n878));
  OR3_X1    g692(.A1(new_n865), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n873), .A2(new_n876), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n860), .A2(KEYINPUT51), .A3(new_n871), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n850), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n313), .A2(new_n765), .A3(new_n394), .A4(new_n517), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n851), .B(KEYINPUT49), .Z(new_n886));
  INV_X1    g700(.A(new_n692), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n680), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n358), .A2(new_n365), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n385), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT55), .Z(new_n892));
  AOI21_X1  g706(.A(new_n847), .B1(new_n838), .B2(new_n839), .ZN(new_n893));
  INV_X1    g707(.A(G210), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n188), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n895), .B2(KEYINPUT56), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n291), .A2(G952), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT123), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT53), .B1(new_n823), .B2(new_n825), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n900), .B(G902), .C1(new_n901), .C2(new_n847), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT122), .B1(new_n893), .B2(new_n188), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n384), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(G51));
  XNOR2_X1  g720(.A(new_n893), .B(KEYINPUT54), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n311), .B(KEYINPUT57), .ZN(new_n908));
  OAI22_X1  g722(.A1(new_n907), .A2(new_n908), .B1(new_n295), .B2(new_n305), .ZN(new_n909));
  INV_X1    g723(.A(new_n782), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n897), .B1(new_n909), .B2(new_n911), .ZN(G54));
  AND2_X1   g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n902), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n915));
  INV_X1    g729(.A(new_n557), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n902), .A2(new_n903), .A3(new_n557), .A4(new_n913), .ZN(new_n919));
  INV_X1    g733(.A(new_n897), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n629), .A2(new_n630), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n898), .B1(new_n907), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n850), .A2(new_n925), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n629), .A2(new_n630), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n849), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n515), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n849), .B(new_n932), .C1(new_n659), .C2(new_n660), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n898), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  INV_X1    g752(.A(G224), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n615), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n835), .B2(G953), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n355), .B(new_n357), .C1(G898), .C2(new_n291), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  NAND2_X1  g757(.A1(new_n424), .A2(new_n400), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n423), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT125), .Z(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n552), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n748), .A2(new_n814), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n693), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  AOI21_X1  g765(.A(new_n774), .B1(new_n635), .B2(new_n644), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n702), .A3(new_n683), .A4(new_n684), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n799), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n951), .A2(new_n793), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n948), .B1(new_n955), .B2(G953), .ZN(new_n956));
  INV_X1    g770(.A(new_n760), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n763), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n702), .A2(new_n815), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n790), .B2(new_n959), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n957), .A2(new_n960), .A3(new_n793), .A4(new_n799), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n291), .ZN(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n947), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n291), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n956), .A2(new_n964), .A3(KEYINPUT126), .A4(new_n966), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G72));
  INV_X1    g785(.A(new_n690), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n441), .A2(new_n408), .A3(new_n416), .ZN(new_n973));
  XOR2_X1   g787(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n842), .A2(new_n843), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n961), .A2(new_n835), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n951), .A2(new_n793), .A3(new_n835), .A4(new_n954), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n972), .B1(new_n981), .B2(new_n976), .ZN(new_n982));
  NOR4_X1   g796(.A1(new_n978), .A2(new_n980), .A3(new_n982), .A4(new_n897), .ZN(G57));
endmodule


