//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G58), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n215), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n250), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n254), .A2(new_n259), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(new_n252), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n263), .A2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n219), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(G58), .A2(G68), .ZN(new_n274));
  OAI21_X1  g0074(.A(G20), .B1(new_n274), .B2(new_n201), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT75), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G159), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n279), .B(G20), .C1(new_n274), .C2(new_n201), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n262), .B1(new_n282), .B2(KEYINPUT16), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT77), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(new_n278), .ZN(new_n285));
  XNOR2_X1  g0085(.A(G58), .B(G68), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n279), .B1(new_n286), .B2(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n270), .A2(new_n215), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT76), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(new_n268), .B2(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n266), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n269), .A3(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n289), .A2(new_n263), .B1(new_n293), .B2(new_n271), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(new_n294), .B2(new_n219), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n271), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n219), .B1(new_n298), .B2(new_n265), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n284), .B(new_n296), .C1(new_n299), .C2(new_n281), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n283), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n296), .B1(new_n299), .B2(new_n281), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n300), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT78), .A3(new_n283), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n261), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n310));
  INV_X1    g0110(.A(G41), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  AOI21_X1  g0112(.A(G1), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G232), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT79), .ZN(new_n316));
  INV_X1    g0116(.A(new_n310), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n317), .A2(G274), .A3(new_n313), .ZN(new_n318));
  OR2_X1    g0118(.A1(G223), .A2(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(G226), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G87), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n321), .A2(new_n270), .B1(new_n266), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n323), .B2(new_n310), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(G179), .A3(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT18), .B1(new_n309), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n261), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n325), .B2(G190), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n270), .B2(new_n215), .ZN(new_n335));
  INV_X1    g0135(.A(new_n271), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n264), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n288), .A3(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n252), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n303), .B(new_n340), .C1(new_n306), .C2(new_n300), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT78), .B1(new_n307), .B2(new_n283), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n331), .B(new_n334), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n328), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n304), .A2(new_n308), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n331), .A4(new_n334), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n330), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G223), .A2(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G222), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n264), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n221), .B2(new_n264), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n317), .B1(new_n357), .B2(KEYINPUT68), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(KEYINPUT68), .B2(new_n357), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n318), .B1(G226), .B2(new_n314), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(G50), .A3(new_n258), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n277), .A2(G150), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n215), .A2(G33), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n255), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(G20), .B2(new_n203), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n364), .B1(G50), .B2(new_n260), .C1(new_n368), .C2(new_n262), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n361), .B2(G169), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n361), .A2(G190), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT71), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT70), .B1(new_n361), .B2(new_n332), .ZN(new_n375));
  OR3_X1    g0175(.A1(new_n361), .A2(KEYINPUT70), .A3(new_n332), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n369), .B(KEYINPUT9), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n233), .A2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n264), .B(new_n382), .C1(G226), .C2(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G97), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT72), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n317), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT73), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n318), .B1(G238), .B2(new_n314), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT13), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n260), .A2(G68), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n394));
  NAND2_X1  g0194(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n253), .A2(G68), .A3(new_n258), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n221), .B2(new_n366), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n252), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT11), .Z(new_n402));
  NOR2_X1   g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n393), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n391), .B2(G169), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n391), .A2(new_n407), .A3(G169), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n362), .C2(new_n391), .ZN(new_n411));
  INV_X1    g0211(.A(new_n403), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n256), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n366), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n252), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n253), .A2(G77), .A3(new_n258), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(G77), .C2(new_n260), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n318), .B1(G244), .B2(new_n314), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n264), .A2(new_n320), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n421), .A2(new_n233), .B1(new_n422), .B2(new_n264), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n264), .A2(G1698), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n220), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n310), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT69), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n419), .B1(new_n429), .B2(G200), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n392), .B2(new_n429), .ZN(new_n431));
  INV_X1    g0231(.A(G169), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n362), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n419), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AND4_X1   g0236(.A1(new_n352), .A2(new_n381), .A3(new_n413), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n270), .A2(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(KEYINPUT4), .A3(G244), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT82), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT4), .B1(new_n438), .B2(G244), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G283), .ZN(new_n442));
  INV_X1    g0242(.A(G250), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n424), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n317), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n447), .A2(G1), .A3(new_n312), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n311), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G274), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(new_n454), .A3(new_n310), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n310), .B1(new_n448), .B2(new_n449), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G257), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G190), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n422), .A2(KEYINPUT6), .A3(G97), .ZN(new_n462));
  XOR2_X1   g0262(.A(G97), .B(G107), .Z(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(KEYINPUT6), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n422), .B2(new_n294), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n252), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n250), .A2(G97), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n253), .B1(G1), .B2(new_n266), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n253), .B(KEYINPUT80), .C1(G1), .C2(new_n266), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT81), .B(new_n469), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n468), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(G200), .B1(new_n446), .B2(new_n459), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n461), .A2(new_n467), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n467), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n460), .A2(new_n362), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n432), .B1(new_n446), .B2(new_n459), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n264), .A2(new_n215), .A3(G68), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n366), .A2(new_n475), .ZN(new_n489));
  AOI21_X1  g0289(.A(G20), .B1(new_n385), .B2(new_n488), .ZN(new_n490));
  NOR3_X1   g0290(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n491));
  OAI221_X1 g0291(.A(new_n487), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n252), .B1(new_n250), .B2(new_n415), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n474), .A2(G87), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  OAI221_X1 g0296(.A(new_n496), .B1(new_n424), .B2(new_n222), .C1(new_n220), .C2(new_n421), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n310), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n312), .A2(G1), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n454), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n317), .B(new_n500), .C1(G250), .C2(new_n499), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G190), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n415), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n474), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n493), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n432), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n509), .B(new_n510), .C1(G179), .C2(new_n502), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n482), .A2(new_n486), .A3(new_n506), .A4(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n442), .B(new_n215), .C1(G33), .C2(new_n475), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n252), .C1(new_n215), .C2(G116), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT20), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n250), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n470), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT85), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n455), .B1(G270), .B2(new_n457), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n264), .A2(G264), .A3(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n264), .A2(G257), .ZN(new_n525));
  OAI221_X1 g0325(.A(new_n523), .B1(new_n524), .B2(new_n264), .C1(new_n525), .C2(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n310), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(G200), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n521), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n432), .B1(new_n522), .B2(new_n527), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n529), .B(G179), .C1(new_n534), .C2(new_n535), .ZN(new_n540));
  INV_X1    g0340(.A(new_n538), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n532), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n264), .A2(new_n215), .A3(G87), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT22), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n215), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n422), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  INV_X1    g0348(.A(new_n496), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n215), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n545), .B2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n252), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n474), .A2(G107), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n250), .A2(new_n422), .ZN(new_n557));
  XOR2_X1   g0357(.A(new_n557), .B(KEYINPUT25), .Z(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n457), .A2(G264), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n525), .A2(new_n320), .B1(new_n266), .B2(new_n561), .ZN(new_n562));
  OR3_X1    g0362(.A1(new_n421), .A2(KEYINPUT87), .A3(new_n443), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT87), .B1(new_n421), .B2(new_n443), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n456), .B(new_n560), .C1(new_n565), .C2(new_n317), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT88), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n566), .A2(new_n567), .A3(new_n362), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n566), .A2(G169), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n566), .B2(new_n362), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n559), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n556), .A2(new_n558), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n551), .B(KEYINPUT24), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(G200), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n566), .A2(new_n392), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n512), .A2(new_n543), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n437), .A2(new_n579), .ZN(G372));
  NAND2_X1  g0380(.A1(new_n379), .A2(new_n380), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n330), .A2(KEYINPUT91), .A3(new_n348), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT91), .B1(new_n330), .B2(new_n348), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n345), .A2(new_n350), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n410), .B1(new_n362), .B2(new_n391), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n412), .B1(new_n587), .B2(new_n408), .ZN(new_n588));
  INV_X1    g0388(.A(new_n435), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n405), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n581), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n371), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n482), .A2(new_n486), .ZN(new_n595));
  INV_X1    g0395(.A(new_n511), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT89), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n495), .A2(new_n597), .A3(new_n505), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n505), .A2(new_n493), .A3(new_n494), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(KEYINPUT89), .B1(G190), .B2(new_n503), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT90), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n595), .A2(new_n601), .A3(new_n602), .A4(new_n577), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n482), .A2(new_n486), .A3(new_n577), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(KEYINPUT89), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n605), .A3(new_n504), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n511), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT90), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n540), .A2(new_n542), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n541), .B1(new_n520), .B2(new_n533), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n571), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(new_n486), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n601), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n506), .A2(new_n511), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT26), .B1(new_n486), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n616), .A2(new_n511), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n437), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n594), .A2(new_n621), .ZN(G369));
  NAND3_X1  g0422(.A1(new_n257), .A2(new_n215), .A3(G13), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n571), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT94), .ZN(new_n630));
  INV_X1    g0430(.A(new_n571), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n628), .ZN(new_n632));
  INV_X1    g0432(.A(new_n628), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT93), .B1(new_n574), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT93), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n559), .A2(new_n635), .A3(new_n628), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n571), .A2(new_n634), .A3(new_n577), .A4(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n630), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n632), .A2(new_n637), .A3(new_n630), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n611), .A2(new_n628), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n629), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n521), .A2(new_n633), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT92), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n543), .B2(new_n645), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(KEYINPUT92), .A3(new_n645), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(G330), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(G399));
  INV_X1    g0451(.A(new_n208), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G41), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(G1), .A2(new_n654), .A3(new_n516), .A4(new_n491), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n213), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT28), .Z(new_n657));
  NAND4_X1  g0457(.A1(new_n612), .A2(new_n595), .A3(new_n577), .A4(new_n601), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n607), .B2(new_n486), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n486), .A2(new_n617), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n596), .B1(new_n660), .B2(new_n614), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(KEYINPUT29), .A3(new_n633), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n628), .B1(new_n613), .B2(new_n619), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(KEYINPUT29), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n528), .A2(new_n362), .A3(new_n502), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n565), .A2(new_n317), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(G264), .B2(new_n457), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n668), .A3(new_n460), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n666), .A2(KEYINPUT30), .A3(new_n668), .A4(new_n460), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n529), .A2(G179), .A3(new_n503), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n566), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n671), .B(new_n672), .C1(new_n460), .C2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT95), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n579), .A2(new_n633), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT95), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n628), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n678), .A2(new_n679), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n665), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n657), .B1(new_n688), .B2(G1), .ZN(G364));
  NOR2_X1   g0489(.A1(new_n249), .A2(G20), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n257), .B1(new_n690), .B2(G45), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n653), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n649), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n648), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n543), .A2(new_n645), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n646), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n249), .A2(new_n266), .A3(KEYINPUT96), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(G13), .B2(G33), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G20), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n693), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n214), .B1(G20), .B2(new_n432), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n215), .A2(G179), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(G190), .A3(G200), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n322), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n215), .A2(new_n362), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G200), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n392), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n714), .B1(G50), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n392), .A3(new_n332), .ZN(new_n719));
  INV_X1    g0519(.A(G159), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT32), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n719), .A2(KEYINPUT32), .A3(new_n720), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n392), .A2(G179), .A3(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n215), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n475), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n712), .A2(new_n392), .A3(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n422), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n716), .A2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n729), .B(new_n264), .C1(new_n219), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G58), .ZN(new_n733));
  INV_X1    g0533(.A(new_n715), .ZN(new_n734));
  AOI21_X1  g0534(.A(G200), .B1(new_n734), .B2(KEYINPUT97), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(KEYINPUT97), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n392), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n736), .A2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n733), .A2(new_n738), .B1(new_n740), .B2(new_n221), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n723), .B(new_n732), .C1(new_n741), .C2(KEYINPUT98), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(KEYINPUT98), .B2(new_n741), .ZN(new_n743));
  INV_X1    g0543(.A(G317), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT33), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n744), .A2(KEYINPUT33), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n730), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G326), .ZN(new_n748));
  INV_X1    g0548(.A(new_n717), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n747), .B1(new_n524), .B2(new_n713), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n725), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n264), .B(new_n750), .C1(G294), .C2(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G311), .A2(new_n739), .B1(new_n737), .B2(G322), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  INV_X1    g0554(.A(G329), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n727), .A2(new_n754), .B1(new_n719), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n752), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n711), .B1(new_n743), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n705), .A2(new_n710), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n208), .A2(G355), .A3(new_n264), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n652), .A2(new_n264), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G45), .B2(new_n212), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n247), .A2(new_n312), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n761), .B1(G116), .B2(new_n208), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n709), .B(new_n759), .C1(new_n760), .C2(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n694), .A2(new_n699), .B1(new_n708), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  INV_X1    g0568(.A(KEYINPUT101), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n589), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n435), .A2(KEYINPUT101), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n419), .A2(new_n628), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT102), .Z(new_n773));
  NAND4_X1  g0573(.A1(new_n770), .A2(new_n431), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n664), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n435), .B2(new_n633), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n664), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n693), .B1(new_n778), .B2(new_n686), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n686), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n704), .A2(new_n711), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n693), .B1(G77), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT100), .ZN(new_n783));
  INV_X1    g0583(.A(new_n719), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n264), .B(new_n726), .C1(G311), .C2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G116), .A2(new_n739), .B1(new_n737), .B2(G294), .ZN(new_n786));
  INV_X1    g0586(.A(new_n713), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n717), .A2(G303), .B1(new_n787), .B2(G107), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n727), .A2(new_n322), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G283), .B2(new_n730), .ZN(new_n790));
  AND4_X1   g0590(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n730), .A2(G150), .B1(new_n717), .B2(G137), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n740), .B2(new_n720), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G143), .B2(new_n737), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT34), .Z(new_n795));
  NOR2_X1   g0595(.A1(new_n727), .A2(new_n219), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n264), .B1(new_n719), .B2(new_n797), .C1(new_n725), .C2(new_n733), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G50), .C2(new_n787), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n791), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n783), .B1(new_n711), .B2(new_n800), .C1(new_n777), .C2(new_n704), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n780), .A2(new_n801), .ZN(G384));
  NOR2_X1   g0602(.A1(new_n690), .A2(new_n257), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n770), .A2(new_n771), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n633), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(KEYINPUT104), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(KEYINPUT104), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n776), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n412), .B(new_n628), .C1(new_n411), .C2(new_n406), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n412), .A2(new_n628), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n588), .A2(new_n405), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n346), .A2(new_n328), .ZN(new_n816));
  INV_X1    g0616(.A(new_n626), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n346), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT37), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n816), .A2(new_n818), .A3(new_n819), .A4(new_n343), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n283), .B1(KEYINPUT16), .B2(new_n282), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n331), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT105), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT105), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(new_n824), .A3(new_n331), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n328), .A2(new_n817), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n343), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n826), .A2(new_n626), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n351), .A2(KEYINPUT106), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT106), .B1(new_n351), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT38), .B(new_n830), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n815), .A2(new_n838), .B1(new_n585), .B2(new_n626), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n330), .A2(new_n348), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n831), .B1(new_n840), .B2(new_n586), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n351), .A2(KEYINPUT106), .A3(new_n831), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT38), .B1(new_n845), .B2(new_n830), .ZN(new_n846));
  INV_X1    g0646(.A(new_n837), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT39), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT39), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n345), .B(new_n350), .C1(new_n582), .C2(new_n583), .ZN(new_n850));
  INV_X1    g0650(.A(new_n818), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n816), .A2(new_n818), .A3(new_n343), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n850), .A2(new_n851), .B1(new_n820), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n849), .B(new_n837), .C1(new_n854), .C2(KEYINPUT38), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n848), .A2(KEYINPUT107), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n411), .A2(new_n412), .A3(new_n633), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT107), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n838), .A2(new_n859), .A3(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n839), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n437), .B(new_n663), .C1(KEYINPUT29), .C2(new_n664), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n594), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n437), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT108), .Z(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n837), .B1(new_n854), .B2(KEYINPUT38), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n813), .A2(new_n866), .A3(new_n777), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n813), .A2(new_n866), .A3(new_n777), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n837), .B2(new_n836), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(G330), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n803), .B1(new_n865), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n865), .B2(new_n878), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n212), .A2(new_n221), .A3(new_n274), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n219), .A2(G50), .ZN(new_n882));
  OAI211_X1 g0682(.A(G1), .B(new_n249), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(G116), .A3(new_n216), .A4(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n880), .A2(new_n883), .A3(new_n888), .ZN(G367));
  INV_X1    g0689(.A(new_n640), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n642), .B1(new_n890), .B2(new_n638), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n483), .A2(new_n628), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n595), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n615), .A2(new_n628), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT42), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n486), .B1(new_n893), .B2(new_n571), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n633), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n891), .A2(KEYINPUT42), .A3(new_n896), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n511), .A2(new_n495), .A3(new_n633), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT109), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n601), .B1(new_n495), .B2(new_n633), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT43), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n902), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n650), .A2(new_n896), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n900), .A2(new_n908), .A3(new_n907), .A4(new_n901), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n653), .B(KEYINPUT41), .Z(new_n917));
  INV_X1    g0717(.A(new_n629), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n891), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT44), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT44), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n921), .B(new_n895), .C1(new_n891), .C2(new_n918), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n919), .B2(new_n896), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n643), .A2(new_n895), .A3(new_n924), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n649), .B(new_n641), .C1(new_n923), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n921), .B1(new_n643), .B2(new_n895), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n919), .A2(KEYINPUT44), .A3(new_n896), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(new_n650), .A3(new_n927), .A4(new_n926), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT111), .ZN(new_n934));
  AND4_X1   g0734(.A1(new_n934), .A2(new_n647), .A3(G330), .A4(new_n648), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n639), .B(new_n640), .C1(new_n611), .C2(new_n628), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n936), .B2(new_n891), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n697), .B2(G330), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(new_n935), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n641), .A2(new_n642), .ZN(new_n940));
  INV_X1    g0740(.A(new_n891), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n937), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n688), .A3(KEYINPUT112), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT112), .ZN(new_n945));
  INV_X1    g0745(.A(new_n935), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n940), .B2(new_n941), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n891), .B(new_n936), .C1(new_n938), .C2(new_n935), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n945), .B1(new_n949), .B2(new_n687), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n929), .A2(new_n933), .A3(new_n944), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n917), .B1(new_n951), .B2(new_n688), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n916), .B1(new_n952), .B2(new_n692), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n240), .A2(new_n652), .A3(new_n264), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n760), .B1(new_n208), .B2(new_n415), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n693), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n270), .B1(new_n719), .B2(new_n744), .C1(new_n731), .C2(new_n561), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n713), .A2(new_n516), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(KEYINPUT46), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT46), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n727), .A2(new_n475), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n725), .A2(new_n422), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(G311), .C2(new_n717), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n738), .B2(new_n524), .C1(new_n754), .C2(new_n740), .ZN(new_n964));
  INV_X1    g0764(.A(G137), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n719), .A2(new_n965), .B1(new_n713), .B2(new_n733), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT113), .Z(new_n967));
  INV_X1    g0767(.A(G150), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(new_n738), .B2(new_n968), .C1(new_n202), .C2(new_n740), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n730), .A2(G159), .B1(new_n717), .B2(G143), .ZN(new_n970));
  INV_X1    g0770(.A(new_n727), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(G77), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n725), .A2(new_n219), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n264), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n960), .A2(new_n964), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n956), .B1(new_n977), .B2(new_n710), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n906), .B2(new_n706), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n953), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT114), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(G387));
  NAND2_X1  g0784(.A1(new_n944), .A2(new_n950), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n985), .B(new_n653), .C1(new_n688), .C2(new_n943), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n943), .A2(new_n692), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n236), .A2(new_n312), .A3(new_n264), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT50), .B1(new_n255), .B2(G50), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n312), .C1(new_n219), .C2(new_n221), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n270), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n516), .A3(new_n491), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n652), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n760), .B1(new_n422), .B2(new_n208), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n693), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G50), .A2(new_n737), .B1(new_n739), .B2(G68), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n270), .B(new_n961), .C1(G150), .C2(new_n784), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n717), .A2(G159), .B1(new_n787), .B2(G77), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n507), .A2(new_n751), .B1(new_n730), .B2(new_n256), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n725), .A2(new_n754), .B1(new_n713), .B2(new_n561), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n730), .A2(G311), .B1(new_n717), .B2(G322), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n738), .B2(new_n744), .C1(new_n524), .C2(new_n740), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT49), .Z(new_n1008));
  OAI221_X1 g0808(.A(new_n270), .B1(new_n719), .B2(new_n748), .C1(new_n516), .C2(new_n727), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n996), .B1(new_n1010), .B2(new_n710), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n641), .B2(new_n706), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n986), .A2(new_n987), .A3(new_n1012), .ZN(G393));
  NAND2_X1  g0813(.A1(new_n929), .A2(new_n933), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n985), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n653), .A3(new_n951), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n929), .A2(new_n933), .A3(new_n692), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n762), .A2(new_n244), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n760), .B1(new_n475), .B2(new_n208), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n693), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n737), .A2(G311), .B1(G317), .B2(new_n717), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n731), .A2(new_n524), .B1(new_n754), .B2(new_n713), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G116), .B2(new_n751), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n264), .B(new_n728), .C1(G322), .C2(new_n784), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n561), .C2(new_n740), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n737), .A2(G159), .B1(G150), .B2(new_n717), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n739), .A2(new_n256), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n270), .B(new_n789), .C1(G143), .C2(new_n784), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n787), .A2(G68), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G77), .A2(new_n751), .B1(new_n730), .B2(G50), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1022), .A2(new_n1026), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1020), .B1(new_n1034), .B2(new_n710), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n895), .B2(new_n706), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1017), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1016), .A2(new_n1037), .ZN(G390));
  AND2_X1   g0838(.A1(new_n813), .A2(new_n777), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n866), .A2(G330), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n858), .B1(new_n808), .B2(new_n813), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n856), .B2(new_n860), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n662), .A2(new_n633), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1045), .A2(new_n775), .B1(new_n633), .B2(new_n804), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n857), .B1(new_n1046), .B2(new_n814), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n870), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1042), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n685), .A2(new_n813), .A3(G330), .A4(new_n777), .ZN(new_n1052));
  AOI211_X1 g0852(.A(KEYINPUT107), .B(new_n849), .C1(new_n836), .C2(new_n837), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n859), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n855), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1051), .B(new_n1052), .C1(new_n1055), .C2(new_n1043), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1040), .A2(new_n437), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n863), .A2(new_n594), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n685), .A2(G330), .A3(new_n777), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n814), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1041), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n808), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n866), .A2(new_n777), .A3(G330), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n814), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1059), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1057), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1050), .A2(new_n1056), .A3(new_n1067), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n653), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1050), .A2(new_n1056), .A3(new_n692), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n693), .B1(new_n256), .B2(new_n781), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G97), .A2(new_n739), .B1(new_n737), .B2(G116), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n264), .B(new_n714), .C1(G294), .C2(new_n784), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n796), .B1(G77), .B2(new_n751), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n730), .A2(G107), .B1(new_n717), .B2(G283), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G159), .A2(new_n751), .B1(new_n717), .B2(G128), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT53), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n713), .A2(new_n968), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1083));
  INV_X1    g0883(.A(G125), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n264), .B1(new_n719), .B2(new_n1084), .C1(new_n202), .C2(new_n727), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT116), .Z(new_n1086));
  OAI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(new_n797), .C2(new_n738), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n739), .A2(new_n1089), .B1(G137), .B2(new_n730), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT115), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1078), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1073), .B1(new_n1092), .B2(new_n710), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT117), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1055), .B2(new_n704), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1072), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1071), .A2(new_n1096), .ZN(G378));
  XNOR2_X1  g0897(.A(new_n1059), .B(KEYINPUT119), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1070), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(G330), .B1(new_n872), .B2(new_n874), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n369), .A2(new_n817), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT55), .Z(new_n1102));
  XNOR2_X1  g0902(.A(new_n381), .B(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(G330), .C1(new_n872), .C2(new_n874), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n862), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n839), .A3(new_n861), .A4(new_n1108), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1099), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n654), .B1(new_n1116), .B2(new_n1099), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1106), .A2(new_n703), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n693), .B1(G50), .B2(new_n781), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n270), .B2(new_n311), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G107), .A2(new_n737), .B1(new_n739), .B2(new_n507), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n311), .B(new_n270), .C1(new_n719), .C2(new_n754), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n973), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n730), .A2(G97), .B1(new_n787), .B2(G77), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n727), .A2(new_n733), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G116), .B2(new_n717), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT58), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1122), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n749), .A2(new_n1084), .B1(new_n968), .B2(new_n725), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n731), .A2(new_n797), .B1(new_n713), .B2(new_n1088), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G128), .C2(new_n737), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n965), .B2(new_n740), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n971), .A2(G159), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1131), .B1(new_n1130), .B2(new_n1129), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1120), .B1(new_n1141), .B2(new_n710), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1112), .A2(new_n692), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1118), .A2(new_n1143), .ZN(G375));
  OAI21_X1  g0944(.A(new_n693), .B1(G68), .B2(new_n781), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n813), .A2(new_n704), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n507), .A2(new_n751), .B1(new_n717), .B2(G294), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n730), .A2(G116), .B1(new_n787), .B2(G97), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n264), .B1(new_n784), .B2(G303), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n972), .A4(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n422), .A2(new_n740), .B1(new_n738), .B2(new_n754), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n965), .A2(new_n738), .B1(new_n740), .B2(new_n968), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G132), .A2(new_n717), .B1(new_n730), .B2(new_n1089), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1127), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n270), .B1(new_n784), .B2(G128), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n751), .A2(G50), .B1(new_n787), .B2(G159), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1150), .A2(new_n1151), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1145), .B(new_n1146), .C1(new_n710), .C2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1039), .A2(new_n1040), .B1(new_n1060), .B2(new_n814), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1066), .B1(new_n1160), .B2(new_n809), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n692), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1162), .B2(KEYINPUT120), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1164), .A3(new_n692), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1161), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1059), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n917), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1068), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(G381));
  OR3_X1    g0971(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G390), .B(G381), .C1(new_n1172), .C2(KEYINPUT121), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n983), .B(new_n1173), .C1(KEYINPUT121), .C2(new_n1172), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT122), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n1112), .A2(new_n692), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1179));
  INV_X1    g0979(.A(G378), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1175), .A2(new_n1181), .ZN(G407));
  NAND2_X1  g0982(.A1(new_n627), .A2(G213), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G213), .B(new_n1184), .C1(new_n1175), .C2(new_n1181), .ZN(G409));
  INV_X1    g0985(.A(G390), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n981), .A2(new_n982), .A3(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n953), .A2(G390), .A3(new_n979), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(G393), .B(new_n767), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n980), .A2(new_n1186), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n953), .A2(G390), .A3(new_n979), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT127), .B1(new_n1194), .B2(new_n1189), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G390), .B1(new_n953), .B2(new_n979), .ZN(new_n1196));
  OAI211_X1 g0996(.A(KEYINPUT127), .B(new_n1189), .C1(new_n1188), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT124), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1099), .A2(new_n1169), .A3(new_n1112), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1143), .A2(new_n1202), .A3(new_n1071), .A4(new_n1096), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1183), .B(new_n1203), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT60), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1168), .B1(new_n1067), .B2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1063), .A2(new_n1059), .A3(KEYINPUT60), .A4(new_n1066), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n653), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(G384), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(KEYINPUT123), .A3(new_n1166), .A4(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1209), .A2(KEYINPUT123), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(KEYINPUT123), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1163), .B1(KEYINPUT120), .B2(new_n1162), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n653), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT60), .B1(new_n1167), .B2(new_n1059), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n1168), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1211), .B(new_n1212), .C1(new_n1213), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1210), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1201), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G375), .A2(G378), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1203), .A2(new_n1183), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(KEYINPUT124), .A4(new_n1218), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT62), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  INV_X1    g1025(.A(G2897), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1183), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1210), .A2(new_n1217), .A3(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n627), .A2(KEYINPUT126), .A3(G213), .A4(G2897), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1227), .B1(new_n1210), .B2(new_n1217), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT61), .B1(new_n1204), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT62), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1200), .B1(new_n1224), .B2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1220), .A2(new_n1223), .A3(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1221), .A2(new_n1222), .A3(KEYINPUT63), .A4(new_n1218), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(new_n1233), .A3(new_n1199), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1240), .ZN(G405));
  NAND2_X1  g1041(.A1(new_n1221), .A2(new_n1181), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1219), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1221), .A2(new_n1181), .A3(new_n1218), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1200), .ZN(G402));
endmodule


