//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT7), .ZN(new_n203));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  INV_X1    g004(.A(G92gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(KEYINPUT8), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G99gat), .B(G106gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  OR2_X1    g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G57gat), .B(G64gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT97), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(KEYINPUT9), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(new_n212), .A3(new_n213), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n211), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n220), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n210), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT10), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n218), .A4(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G230gat), .ZN(new_n228));
  INV_X1    g027(.A(G233gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n221), .A2(new_n223), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  XNOR2_X1  g033(.A(G120gat), .B(G148gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G176gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G204gat), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT101), .ZN(new_n242));
  INV_X1    g041(.A(G29gat), .ZN(new_n243));
  INV_X1    g042(.A(G36gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT14), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G29gat), .B2(G36gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT14), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248));
  INV_X1    g047(.A(G50gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G43gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n250), .B2(KEYINPUT90), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G43gat), .B(G50gat), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n246), .A2(new_n247), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n252), .B(new_n253), .C1(new_n254), .C2(KEYINPUT15), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n252), .A2(new_n253), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n210), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT41), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT100), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n211), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT100), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT91), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n210), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n266), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n266), .B2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(G218gat), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n266), .A2(new_n274), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G190gat), .ZN(new_n282));
  AOI21_X1  g081(.A(G218gat), .B1(new_n282), .B2(new_n276), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n242), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n279), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(G218gat), .A3(new_n276), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT101), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT99), .B(G134gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G162gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n258), .A2(KEYINPUT41), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT101), .A4(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT21), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n222), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT16), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(G1gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G1gat), .B2(new_n302), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(G8gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n222), .B2(new_n297), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT98), .B(G155gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n301), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n312));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n311), .B(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n296), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n279), .ZN(new_n319));
  NAND2_X1  g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n322));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n320), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n321), .B(new_n323), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(KEYINPUT74), .A3(new_n321), .A4(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n317), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  INV_X1    g136(.A(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G141gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(G141gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n336), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G155gat), .B(G162gat), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT2), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n348), .B2(KEYINPUT2), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT77), .B(G141gat), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT78), .B(new_n343), .C1(new_n354), .C2(new_n337), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n345), .A2(new_n347), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n338), .A2(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n358), .A3(KEYINPUT76), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n349), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n346), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n357), .B1(new_n356), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n335), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n356), .A2(new_n317), .A3(new_n364), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n334), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n356), .B2(new_n364), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n356), .A2(new_n375), .A3(new_n364), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n335), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  OAI21_X1  g179(.A(G22gat), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n382));
  INV_X1    g181(.A(G22gat), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n356), .A2(new_n375), .A3(new_n364), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n376), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n385), .A2(new_n335), .B1(new_n334), .B2(new_n372), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n382), .B(new_n383), .C1(new_n386), .C2(new_n369), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(KEYINPUT87), .A3(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G78gat), .B(G106gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT31), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(new_n249), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n380), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n383), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n381), .A2(KEYINPUT86), .A3(new_n387), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n397), .A3(new_n383), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT85), .ZN(new_n401));
  INV_X1    g200(.A(new_n391), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n395), .A2(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT75), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G64gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(new_n206), .ZN(new_n407));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT68), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410));
  AND2_X1   g209(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414));
  INV_X1    g213(.A(G183gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n418), .A3(new_n275), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT28), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT28), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n275), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n409), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g224(.A(KEYINPUT68), .B(new_n423), .C1(new_n419), .C2(KEYINPUT28), .ZN(new_n426));
  NOR2_X1   g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT26), .ZN(new_n428));
  NAND2_X1  g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT65), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n425), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n427), .B(KEYINPUT23), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n430), .A2(new_n436), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n432), .B(KEYINPUT24), .ZN(new_n441));
  NOR2_X1   g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n435), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n442), .B(KEYINPUT64), .Z(new_n446));
  INV_X1    g245(.A(new_n441), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n445), .B(new_n430), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n439), .A2(new_n444), .B1(new_n448), .B2(new_n440), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n371), .B(new_n408), .C1(new_n434), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n334), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n420), .A2(new_n424), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT68), .ZN(new_n453));
  INV_X1    g252(.A(new_n433), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n420), .A2(new_n409), .A3(new_n424), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n438), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n445), .A3(new_n444), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n440), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n456), .A2(new_n460), .A3(G226gat), .A4(G233gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(new_n451), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n451), .B1(new_n450), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n407), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  INV_X1    g265(.A(new_n407), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n468), .A3(KEYINPUT30), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n407), .C1(new_n463), .C2(new_n464), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT72), .ZN(new_n473));
  XNOR2_X1  g272(.A(G113gat), .B(G120gat), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT69), .B(G127gat), .C1(new_n474), .C2(KEYINPUT1), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT1), .ZN(new_n476));
  INV_X1    g275(.A(G127gat), .ZN(new_n477));
  INV_X1    g276(.A(G113gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(G120gat), .ZN(new_n479));
  INV_X1    g278(.A(G120gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(G113gat), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n476), .B(new_n477), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G134gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n475), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n475), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n434), .B2(new_n449), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n456), .A2(new_n460), .A3(new_n486), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(G227gat), .A2(G233gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n473), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT34), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n473), .B(new_n494), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n491), .A3(new_n489), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n488), .A2(KEYINPUT70), .A3(new_n489), .A4(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT33), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G43gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G71gat), .ZN(new_n506));
  INV_X1    g305(.A(G99gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(KEYINPUT33), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT32), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n510), .B(new_n512), .C1(new_n499), .C2(new_n500), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n501), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n510), .ZN(new_n517));
  AND4_X1   g316(.A1(new_n496), .A2(new_n509), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT71), .B1(new_n501), .B2(new_n515), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n513), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n496), .B1(new_n520), .B2(new_n509), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n403), .B(new_n472), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n487), .B1(new_n384), .B2(new_n376), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n356), .A2(new_n364), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n486), .A2(new_n526), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT3), .B1(new_n366), .B2(new_n367), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n486), .A3(new_n370), .ZN(new_n530));
  NAND2_X1  g329(.A1(G225gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n367), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n317), .B1(new_n535), .B2(new_n365), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n370), .A2(new_n486), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n365), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n527), .B1(new_n541), .B2(new_n486), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n532), .B1(new_n542), .B2(new_n531), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n534), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G85gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT6), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n534), .C1(new_n540), .C2(new_n543), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n544), .A2(KEYINPUT6), .A3(new_n550), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT35), .B1(new_n522), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n382), .B1(new_n386), .B2(new_n369), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n393), .B1(new_n558), .B2(G22gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n402), .B1(new_n559), .B2(new_n387), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n400), .A2(new_n560), .A3(new_n394), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n401), .A2(new_n402), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n514), .A2(new_n509), .A3(new_n517), .ZN(new_n564));
  INV_X1    g363(.A(new_n496), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n520), .A2(new_n496), .A3(new_n509), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n551), .A2(KEYINPUT88), .A3(new_n552), .A4(new_n553), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n555), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n472), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n472), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n542), .A2(new_n531), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n528), .A2(new_n530), .ZN(new_n578));
  OAI211_X1 g377(.A(KEYINPUT39), .B(new_n577), .C1(new_n578), .C2(new_n531), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n531), .B1(new_n528), .B2(new_n530), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n549), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n579), .A2(KEYINPUT40), .A3(new_n549), .A4(new_n582), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n576), .A2(new_n551), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n463), .B2(new_n464), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n466), .A2(KEYINPUT37), .A3(new_n462), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n467), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT38), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .A4(new_n467), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n465), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n587), .B(new_n403), .C1(new_n573), .C2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n563), .B1(new_n556), .B2(new_n576), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n566), .A2(KEYINPUT36), .A3(new_n567), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n518), .B2(new_n521), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n273), .A2(new_n307), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n262), .A2(new_n306), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n262), .A2(new_n306), .A3(KEYINPUT92), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(KEYINPUT93), .B(KEYINPUT18), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n273), .A2(new_n307), .B1(new_n606), .B2(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G197gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT11), .ZN(new_n619));
  INV_X1    g418(.A(G169gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  NOR2_X1   g421(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n262), .B2(new_n306), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n307), .A2(KEYINPUT94), .A3(new_n255), .A4(new_n256), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n610), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n616), .A2(KEYINPUT95), .A3(new_n622), .A4(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n614), .B1(new_n613), .B2(new_n610), .ZN(new_n632));
  AND4_X1   g431(.A1(new_n610), .A2(new_n603), .A3(new_n608), .A4(new_n614), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n630), .B(new_n622), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n616), .A2(new_n630), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n622), .B(KEYINPUT89), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT96), .B1(new_n602), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n643), .B(new_n644), .C1(new_n575), .C2(new_n601), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n241), .B(new_n316), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n556), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n576), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  AND2_X1   g450(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n656), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n650), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n656), .B2(KEYINPUT42), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(G1325gat));
  INV_X1    g459(.A(G15gat), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n600), .A2(new_n598), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n646), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n518), .A2(new_n521), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n661), .B2(new_n666), .ZN(G1326gat));
  INV_X1    g466(.A(new_n316), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n602), .A2(new_n641), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n643), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n602), .A2(KEYINPUT96), .A3(new_n641), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n241), .A4(new_n563), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n646), .B2(new_n403), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT43), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n677), .A2(G22gat), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(G22gat), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(G1327gat));
  AOI21_X1  g481(.A(KEYINPUT106), .B1(new_n293), .B2(new_n294), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n293), .A2(KEYINPUT106), .A3(new_n294), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n575), .A2(KEYINPUT105), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n557), .A2(new_n574), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n601), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n662), .A2(KEYINPUT104), .A3(new_n597), .A4(new_n596), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n688), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n687), .B1(new_n602), .B2(new_n296), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n315), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n240), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n641), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n556), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n670), .A2(new_n671), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n296), .A3(new_n701), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n243), .A3(new_n556), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n706), .A2(G36gat), .A3(new_n472), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n702), .B2(new_n472), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(G1329gat));
  OAI21_X1  g516(.A(G43gat), .B1(new_n702), .B2(new_n662), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n707), .A2(new_n719), .A3(new_n665), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT47), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1330gat));
  OAI21_X1  g525(.A(G50gat), .B1(new_n702), .B2(new_n403), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n707), .A2(new_n249), .A3(new_n563), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  AOI22_X1  g531(.A1(new_n689), .A2(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n316), .A2(new_n644), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n556), .B(KEYINPUT108), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n240), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n735), .B2(new_n240), .ZN(new_n740));
  NOR4_X1   g539(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT109), .A4(new_n241), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n576), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n742), .A2(new_n576), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g546(.A1(new_n735), .A2(new_n240), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(G71gat), .A3(new_n664), .ZN(new_n749));
  INV_X1    g548(.A(new_n662), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n740), .B2(new_n741), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(G71gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n563), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT110), .B(G78gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n697), .A2(new_n698), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n700), .A2(new_n641), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n240), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n703), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n601), .A2(new_n693), .ZN(new_n764));
  INV_X1    g563(.A(new_n695), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n557), .A2(new_n690), .A3(new_n574), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n690), .B1(new_n557), .B2(new_n574), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n758), .A2(new_n296), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n763), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n763), .B(new_n772), .C1(new_n733), .C2(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n769), .B1(new_n692), .B2(new_n696), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(KEYINPUT51), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n733), .A2(KEYINPUT111), .A3(new_n772), .A4(new_n769), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n773), .A2(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n205), .A3(new_n556), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n762), .B1(new_n781), .B2(new_n241), .ZN(G1336gat));
  INV_X1    g581(.A(new_n759), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n576), .B(new_n783), .C1(new_n697), .C2(new_n698), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n777), .B(new_n772), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n576), .A2(new_n206), .A3(new_n240), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT113), .Z(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  INV_X1    g590(.A(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n780), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n784), .B2(G92gat), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n777), .A2(new_n776), .A3(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT112), .B1(new_n777), .B2(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n774), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n788), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n790), .B1(new_n795), .B2(new_n805), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n761), .B2(new_n662), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n780), .A2(new_n507), .A3(new_n665), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n241), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n403), .A2(G106gat), .A3(new_n241), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n786), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n760), .B2(new_n563), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n780), .A2(new_n810), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(G1339gat));
  NOR2_X1   g618(.A1(new_n734), .A2(new_n240), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n627), .A2(new_n629), .B1(new_n613), .B2(new_n610), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n621), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n637), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n232), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n827));
  NAND3_X1  g626(.A1(new_n227), .A2(new_n231), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(KEYINPUT117), .A3(new_n237), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT117), .B1(new_n828), .B2(new_n237), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT55), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n238), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n293), .A2(KEYINPUT106), .A3(new_n294), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n683), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n836), .B(new_n840), .C1(new_n837), .C2(new_n683), .ZN(new_n841));
  INV_X1    g640(.A(new_n686), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n644), .A2(new_n835), .B1(new_n241), .B2(new_n824), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n839), .A2(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n821), .B1(new_n844), .B2(new_n700), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n568), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n703), .A2(new_n576), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n644), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n845), .A2(new_n736), .ZN(new_n850));
  INV_X1    g649(.A(new_n522), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n478), .A3(new_n851), .A4(new_n641), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT119), .ZN(G1340gat));
  AND2_X1   g653(.A1(new_n850), .A2(new_n851), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n480), .A3(new_n240), .ZN(new_n856));
  OAI21_X1  g655(.A(G120gat), .B1(new_n848), .B2(new_n241), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n855), .B2(new_n700), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n848), .A2(new_n477), .A3(new_n315), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(G1342gat));
  NOR2_X1   g660(.A1(new_n295), .A2(new_n576), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n845), .A2(new_n736), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT69), .B(G134gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n568), .A4(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n568), .A3(new_n736), .A4(new_n863), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT121), .B1(new_n869), .B2(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n848), .B2(new_n295), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n868), .A2(new_n874), .A3(new_n870), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n872), .B(new_n873), .C1(new_n876), .C2(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n843), .A2(new_n295), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n840), .B1(new_n686), .B2(new_n836), .ZN(new_n880));
  INV_X1    g679(.A(new_n841), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n820), .B1(new_n882), .B2(new_n315), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT57), .B1(new_n883), .B2(new_n403), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n845), .A2(new_n885), .A3(new_n563), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n662), .A2(new_n847), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n641), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT123), .B1(new_n888), .B2(new_n354), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n750), .A2(new_n403), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n845), .A2(new_n472), .A3(new_n736), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n641), .A2(new_n338), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n888), .B2(new_n354), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n889), .A2(new_n894), .A3(KEYINPUT58), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  AOI221_X4 g695(.A(new_n893), .B1(KEYINPUT123), .B2(new_n896), .C1(new_n888), .C2(new_n354), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(G1344gat));
  OR2_X1    g697(.A1(new_n891), .A2(G148gat), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n899), .A2(KEYINPUT124), .A3(new_n241), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n899), .B2(new_n241), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n845), .A2(new_n563), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n836), .A2(new_n296), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n700), .B1(new_n879), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n885), .B(new_n563), .C1(new_n907), .C2(new_n820), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n905), .A2(new_n240), .A3(new_n887), .A4(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n887), .A3(new_n886), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n911), .B2(new_n241), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n337), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n902), .B1(new_n910), .B2(new_n913), .ZN(G1345gat));
  INV_X1    g713(.A(G155gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n911), .A2(new_n915), .A3(new_n315), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n891), .A2(new_n315), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(G1346gat));
  OAI21_X1  g717(.A(G162gat), .B1(new_n911), .B2(new_n842), .ZN(new_n919));
  INV_X1    g718(.A(G162gat), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n850), .A2(new_n920), .A3(new_n863), .A4(new_n890), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n736), .A2(new_n472), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n846), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(G169gat), .A3(new_n641), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n845), .A2(new_n703), .A3(new_n568), .A4(new_n576), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n620), .B1(new_n926), .B2(new_n644), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n925), .A2(KEYINPUT125), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT125), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1348gat));
  INV_X1    g729(.A(new_n926), .ZN(new_n931));
  AOI21_X1  g730(.A(G176gat), .B1(new_n931), .B2(new_n240), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n240), .A2(G176gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n924), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n846), .A2(new_n700), .A3(new_n923), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G183gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n413), .A2(new_n418), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(new_n700), .ZN(new_n940));
  NOR4_X1   g739(.A1(new_n926), .A2(KEYINPUT126), .A3(new_n938), .A4(new_n315), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n936), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n275), .A3(new_n686), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n924), .A2(new_n296), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(G190gat), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT61), .B(new_n275), .C1(new_n924), .C2(new_n296), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NAND4_X1  g751(.A1(new_n845), .A2(new_n703), .A3(new_n576), .A4(new_n890), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n641), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n923), .A2(new_n662), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n905), .A2(new_n908), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(new_n641), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n960), .B2(new_n955), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n905), .A2(new_n240), .A3(new_n908), .ZN(new_n962));
  OAI21_X1  g761(.A(G204gat), .B1(new_n962), .B2(new_n957), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n953), .A2(G204gat), .A3(new_n241), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(new_n964), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(new_n964), .ZN(new_n968));
  OAI221_X1 g767(.A(new_n963), .B1(new_n964), .B2(new_n965), .C1(new_n967), .C2(new_n968), .ZN(G1353gat));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n318), .A3(new_n700), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n905), .A2(new_n700), .A3(new_n908), .A4(new_n958), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n954), .B2(new_n686), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n295), .A2(new_n279), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n959), .B2(new_n976), .ZN(G1355gat));
endmodule


