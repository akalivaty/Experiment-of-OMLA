

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594;

  XOR2_X1 U327 ( .A(n470), .B(KEYINPUT28), .Z(n538) );
  XOR2_X1 U328 ( .A(n453), .B(n452), .Z(n535) );
  XOR2_X1 U329 ( .A(n310), .B(n435), .Z(n532) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U331 ( .A(n341), .B(KEYINPUT7), .Z(n296) );
  AND2_X1 U332 ( .A1(n416), .A2(n415), .ZN(n297) );
  INV_X1 U333 ( .A(n530), .ZN(n415) );
  INV_X1 U334 ( .A(KEYINPUT33), .ZN(n320) );
  XNOR2_X1 U335 ( .A(n353), .B(n295), .ZN(n300) );
  XNOR2_X1 U336 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U337 ( .A(n429), .B(n300), .ZN(n304) );
  XNOR2_X1 U338 ( .A(n323), .B(n322), .ZN(n327) );
  NOR2_X1 U339 ( .A1(n538), .A2(n469), .ZN(n544) );
  NOR2_X1 U340 ( .A1(n454), .A2(n546), .ZN(n455) );
  XOR2_X1 U341 ( .A(n583), .B(KEYINPUT41), .Z(n564) );
  INV_X1 U342 ( .A(G29GAT), .ZN(n483) );
  XNOR2_X1 U343 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n488) );
  XNOR2_X1 U344 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U345 ( .A(n489), .B(n488), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U347 ( .A(G211GAT), .B(KEYINPUT21), .Z(n299) );
  XNOR2_X1 U348 ( .A(G197GAT), .B(KEYINPUT84), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n429) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G218GAT), .Z(n353) );
  XOR2_X1 U351 ( .A(KEYINPUT90), .B(G92GAT), .Z(n302) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n306) );
  XOR2_X1 U355 ( .A(G169GAT), .B(G8GAT), .Z(n334) );
  XOR2_X1 U356 ( .A(G176GAT), .B(G64GAT), .Z(n328) );
  XNOR2_X1 U357 ( .A(n334), .B(n328), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n308) );
  XNOR2_X1 U360 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U362 ( .A(KEYINPUT18), .B(n309), .ZN(n435) );
  INV_X1 U363 ( .A(n532), .ZN(n463) );
  XNOR2_X1 U364 ( .A(KEYINPUT67), .B(G204GAT), .ZN(n316) );
  INV_X1 U365 ( .A(G148GAT), .ZN(n311) );
  NAND2_X1 U366 ( .A1(G78GAT), .A2(n311), .ZN(n314) );
  INV_X1 U367 ( .A(G78GAT), .ZN(n312) );
  NAND2_X1 U368 ( .A1(n312), .A2(G148GAT), .ZN(n313) );
  NAND2_X1 U369 ( .A1(n314), .A2(n313), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n427) );
  XOR2_X1 U371 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XNOR2_X1 U372 ( .A(n427), .B(n445), .ZN(n318) );
  AND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n319), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U377 ( .A(n350), .B(KEYINPUT69), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT31), .B(KEYINPUT68), .Z(n325) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(KEYINPUT32), .ZN(n324) );
  XOR2_X1 U380 ( .A(n325), .B(n324), .Z(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n330) );
  XOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT13), .Z(n367) );
  XNOR2_X1 U383 ( .A(n328), .B(n367), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n583) );
  XOR2_X1 U385 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n332) );
  NAND2_X1 U386 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U388 ( .A(n333), .B(KEYINPUT65), .Z(n336) );
  XOR2_X1 U389 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XNOR2_X1 U390 ( .A(n420), .B(n334), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U392 ( .A(G15GAT), .B(G1GAT), .Z(n368) );
  XOR2_X1 U393 ( .A(n337), .B(n368), .Z(n339) );
  XNOR2_X1 U394 ( .A(G113GAT), .B(G197GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n343) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n340), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(G43GAT), .B(G50GAT), .ZN(n342) );
  XOR2_X1 U399 ( .A(n296), .B(n342), .Z(n358) );
  XNOR2_X1 U400 ( .A(n343), .B(n358), .ZN(n578) );
  NAND2_X1 U401 ( .A1(n564), .A2(n578), .ZN(n346) );
  XOR2_X1 U402 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT112), .B(n344), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n381) );
  XOR2_X1 U405 ( .A(KEYINPUT9), .B(KEYINPUT70), .Z(n352) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n348) );
  XNOR2_X1 U407 ( .A(KEYINPUT72), .B(KEYINPUT64), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U411 ( .A(G134GAT), .B(KEYINPUT71), .Z(n406) );
  XOR2_X1 U412 ( .A(n353), .B(n406), .Z(n355) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n360) );
  XOR2_X1 U416 ( .A(G162GAT), .B(G106GAT), .Z(n419) );
  XOR2_X1 U417 ( .A(n358), .B(n419), .Z(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n570) );
  XOR2_X1 U419 ( .A(G211GAT), .B(G71GAT), .Z(n362) );
  XNOR2_X1 U420 ( .A(G183GAT), .B(G127GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n364) );
  XNOR2_X1 U423 ( .A(G64GAT), .B(KEYINPUT75), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U425 ( .A(n366), .B(n365), .Z(n370) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n372) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U432 ( .A(G78GAT), .B(G155GAT), .Z(n376) );
  XNOR2_X1 U433 ( .A(G22GAT), .B(G8GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n377), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n586) );
  INV_X1 U437 ( .A(n586), .ZN(n490) );
  AND2_X1 U438 ( .A1(n570), .A2(n490), .ZN(n380) );
  AND2_X1 U439 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n382), .B(KEYINPUT47), .ZN(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT73), .B(n570), .ZN(n487) );
  XOR2_X1 U442 ( .A(KEYINPUT36), .B(n487), .Z(n591) );
  NOR2_X1 U443 ( .A1(n591), .A2(n490), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT45), .B(n383), .Z(n384) );
  NOR2_X1 U445 ( .A1(n583), .A2(n384), .ZN(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT66), .B(n578), .ZN(n572) );
  INV_X1 U447 ( .A(n572), .ZN(n462) );
  NAND2_X1 U448 ( .A1(n385), .A2(n462), .ZN(n386) );
  NAND2_X1 U449 ( .A1(n387), .A2(n386), .ZN(n389) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n543) );
  NOR2_X1 U452 ( .A1(n463), .A2(n543), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n390), .B(KEYINPUT54), .ZN(n416) );
  XOR2_X1 U454 ( .A(G127GAT), .B(KEYINPUT0), .Z(n392) );
  XNOR2_X1 U455 ( .A(G113GAT), .B(KEYINPUT77), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n444) );
  XOR2_X1 U457 ( .A(n444), .B(KEYINPUT5), .Z(n394) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n414) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n396) );
  XNOR2_X1 U461 ( .A(KEYINPUT89), .B(KEYINPUT87), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U463 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n398) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U466 ( .A(n400), .B(n399), .Z(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n402) );
  XNOR2_X1 U468 ( .A(KEYINPUT85), .B(G155GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U470 ( .A(KEYINPUT2), .B(n403), .Z(n430) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G162GAT), .Z(n405) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(G148GAT), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U474 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G120GAT), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n430), .B(n410), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U479 ( .A(n414), .B(n413), .Z(n530) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n418) );
  XNOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U483 ( .A(G218GAT), .B(n419), .Z(n422) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U486 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U489 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n470) );
  NAND2_X1 U492 ( .A1(n297), .A2(n470), .ZN(n434) );
  XOR2_X1 U493 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n454) );
  INV_X1 U495 ( .A(n435), .ZN(n453) );
  XOR2_X1 U496 ( .A(G190GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G99GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT78), .Z(n439) );
  XNOR2_X1 U500 ( .A(G169GAT), .B(G15GAT), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(KEYINPUT79), .Z(n443) );
  XNOR2_X1 U504 ( .A(KEYINPUT80), .B(KEYINPUT20), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n449) );
  XOR2_X1 U506 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U511 ( .A(n535), .ZN(n546) );
  XOR2_X1 U512 ( .A(KEYINPUT119), .B(n455), .Z(n573) );
  NAND2_X1 U513 ( .A1(n573), .A2(n586), .ZN(n457) );
  XNOR2_X1 U514 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(G1350GAT) );
  NAND2_X1 U516 ( .A1(n573), .A2(n564), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n459) );
  XOR2_X1 U518 ( .A(G176GAT), .B(KEYINPUT56), .Z(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U521 ( .A(KEYINPUT38), .B(KEYINPUT100), .Z(n482) );
  NOR2_X1 U522 ( .A1(n462), .A2(n583), .ZN(n494) );
  XOR2_X1 U523 ( .A(n463), .B(KEYINPUT91), .Z(n464) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n464), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n544), .A2(n546), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n415), .A2(n465), .ZN(n466) );
  XOR2_X1 U527 ( .A(n466), .B(KEYINPUT92), .Z(n476) );
  NAND2_X1 U528 ( .A1(n535), .A2(n532), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n470), .A2(n467), .ZN(n468) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(n468), .Z(n473) );
  INV_X1 U531 ( .A(n469), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n470), .A2(n535), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U534 ( .A1(n472), .A2(n576), .ZN(n559) );
  NAND2_X1 U535 ( .A1(n473), .A2(n559), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n415), .A2(n474), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n476), .A2(n475), .ZN(n493) );
  NAND2_X1 U538 ( .A1(n493), .A2(n490), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT98), .B(n477), .ZN(n478) );
  NOR2_X1 U540 ( .A1(n591), .A2(n478), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT99), .B(KEYINPUT37), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n527) );
  NAND2_X1 U543 ( .A1(n494), .A2(n527), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n511) );
  NAND2_X1 U545 ( .A1(n511), .A2(n530), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT97), .B(KEYINPUT39), .Z(n484) );
  NAND2_X1 U547 ( .A1(n487), .A2(n573), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n497) );
  OR2_X1 U549 ( .A1(n487), .A2(n490), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT16), .B(n491), .Z(n492) );
  AND2_X1 U551 ( .A1(n493), .A2(n492), .ZN(n515) );
  NAND2_X1 U552 ( .A1(n494), .A2(n515), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT93), .B(n495), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n530), .A2(n504), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U556 ( .A1(n532), .A2(n504), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n500) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT94), .B(n501), .Z(n503) );
  NAND2_X1 U562 ( .A1(n504), .A2(n535), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n538), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U566 ( .A1(n532), .A2(n511), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n510) );
  XOR2_X1 U569 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n508) );
  NAND2_X1 U570 ( .A1(n511), .A2(n535), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1330GAT) );
  XOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT103), .Z(n513) );
  NAND2_X1 U574 ( .A1(n511), .A2(n538), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n518) );
  INV_X1 U577 ( .A(n564), .ZN(n514) );
  NOR2_X1 U578 ( .A1(n578), .A2(n514), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n515), .A2(n528), .ZN(n516) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(n516), .Z(n524) );
  NAND2_X1 U581 ( .A1(n530), .A2(n524), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n524), .A2(n532), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(KEYINPUT106), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  XOR2_X1 U587 ( .A(G71GAT), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U588 ( .A1(n535), .A2(n524), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U591 ( .A1(n538), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT108), .B(n529), .Z(n537) );
  NAND2_X1 U595 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n531), .ZN(G1336GAT) );
  XOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT109), .Z(n534) );
  NAND2_X1 U598 ( .A1(n537), .A2(n532), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1339GAT) );
  NOR2_X1 U607 ( .A1(n415), .A2(n543), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n544), .A2(n557), .ZN(n545) );
  NOR2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n572), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(n547), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n549) );
  NAND2_X1 U613 ( .A1(n553), .A2(n564), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G120GAT), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U616 ( .A1(n553), .A2(n586), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n487), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(G134GAT), .B(n556), .Z(G1343GAT) );
  INV_X1 U623 ( .A(n557), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n578), .A2(n568), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n562) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT52), .B(n563), .Z(n566) );
  NAND2_X1 U631 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n586), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U635 ( .A(n568), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(G162GAT), .B(n571), .Z(G1347GAT) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1348GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n297), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT123), .ZN(n589) );
  NAND2_X1 U643 ( .A1(n589), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n589), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .Z(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n589), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(G218GAT), .B(n594), .Z(G1355GAT) );
endmodule

