//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G101), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI211_X1 g009(.A(KEYINPUT78), .B(new_n188), .C1(new_n190), .C2(new_n192), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n188), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n189), .A3(G104), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n191), .A2(KEYINPUT77), .A3(G107), .ZN(new_n201));
  OAI211_X1 g015(.A(KEYINPUT3), .B(new_n200), .C1(new_n201), .C2(new_n199), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT76), .B(new_n203), .C1(new_n190), .C2(KEYINPUT77), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT80), .B1(new_n197), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n191), .A2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n199), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n198), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n189), .A2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n207), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n193), .A2(new_n194), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n225), .B2(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n225), .C2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(G128), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n226), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n206), .A2(new_n220), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n215), .B1(new_n202), .B2(new_n204), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n213), .B(KEYINPUT4), .C1(new_n239), .C2(new_n188), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT0), .A4(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n211), .A2(new_n192), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n188), .A2(KEYINPUT4), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G137), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(G134), .B2(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n250), .A2(KEYINPUT11), .A3(G137), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n229), .A2(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n234), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n227), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n222), .A2(new_n224), .A3(new_n226), .A4(KEYINPUT79), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n213), .A2(new_n219), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n236), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n238), .A2(new_n249), .A3(new_n261), .A4(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n235), .B1(new_n197), .B2(new_n205), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n272), .A2(KEYINPUT12), .A3(new_n260), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT12), .B1(new_n272), .B2(new_n260), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(G227), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n238), .A2(new_n249), .A3(new_n269), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n260), .ZN(new_n282));
  INV_X1    g096(.A(new_n279), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n270), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n187), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n240), .A2(new_n248), .B1(new_n268), .B2(new_n236), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n261), .B1(new_n289), .B2(new_n238), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n273), .A2(new_n274), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n270), .A2(new_n283), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n291), .A2(KEYINPUT82), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n283), .B1(new_n282), .B2(new_n270), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT81), .B(G469), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT83), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(KEYINPUT2), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(KEYINPUT2), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT2), .B(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n313), .A2(new_n320), .A3(KEYINPUT66), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n246), .A2(new_n247), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n188), .B1(new_n211), .B2(new_n192), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n318), .A2(new_n319), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n315), .B2(KEYINPUT5), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(new_n314), .A3(KEYINPUT84), .A4(G116), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n310), .B1(new_n309), .B2(KEYINPUT5), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n206), .A2(new_n220), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g152(.A(G110), .B(G122), .Z(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT85), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n328), .A2(new_n337), .A3(new_n344), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(KEYINPUT6), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n328), .B2(new_n337), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n338), .A2(new_n352), .A3(new_n345), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n348), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT73), .B(G125), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n245), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n232), .A2(G128), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT65), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n234), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n227), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n359), .B1(new_n363), .B2(new_n358), .ZN(new_n364));
  INV_X1    g178(.A(G224), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n364), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n336), .B1(new_n197), .B2(new_n205), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT5), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n331), .A2(new_n372), .A3(G113), .A4(new_n333), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n313), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n213), .A2(new_n374), .A3(new_n219), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n340), .A2(KEYINPUT8), .A3(new_n343), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT8), .B1(new_n340), .B2(new_n343), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n364), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n364), .A2(new_n366), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n235), .A2(new_n357), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(new_n359), .A3(KEYINPUT7), .A4(new_n367), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(KEYINPUT87), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n347), .B1(new_n385), .B2(KEYINPUT87), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n286), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT88), .B(new_n286), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n370), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G210), .B1(G237), .B2(G902), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n370), .A2(new_n390), .A3(new_n393), .A4(new_n391), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n308), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n270), .A2(new_n283), .ZN(new_n398));
  OAI22_X1  g212(.A1(new_n296), .A2(new_n297), .B1(new_n292), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n291), .A2(KEYINPUT82), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n286), .B(new_n301), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n280), .A2(new_n284), .ZN(new_n402));
  OAI21_X1  g216(.A(G469), .B1(new_n402), .B2(G902), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n305), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n306), .A2(new_n397), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(G119), .B(G128), .Z(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT24), .B(G110), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT23), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n314), .B2(G128), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n412), .B(new_n413), .C1(G119), .C2(new_n221), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(G110), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n357), .A2(G140), .ZN(new_n417));
  INV_X1    g231(.A(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G125), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT72), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(KEYINPUT72), .A3(G125), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n223), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(G146), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n416), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(G125), .B(G140), .Z(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G146), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n414), .A2(G110), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n408), .A2(new_n409), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n427), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT74), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G137), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n429), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  INV_X1    g255(.A(new_n435), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n428), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n443), .A3(new_n286), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n440), .A2(new_n443), .A3(KEYINPUT25), .A4(new_n286), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT75), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(G217), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(G234), .B2(new_n286), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n443), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n453), .A2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n449), .A2(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT64), .B1(new_n253), .B2(G134), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT64), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n250), .A3(G137), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n253), .A2(G134), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G131), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n259), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n235), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n245), .B1(new_n259), .B2(new_n257), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n324), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n245), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n260), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n465), .A2(new_n259), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n363), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n321), .A2(new_n323), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n459), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT69), .B1(new_n477), .B2(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT28), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n277), .A3(G210), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT68), .Z(new_n487));
  XNOR2_X1  g301(.A(new_n484), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n479), .A2(new_n481), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT70), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n467), .A2(new_n324), .A3(new_n468), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n474), .B1(new_n471), .B2(new_n473), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT28), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n488), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT30), .B1(new_n467), .B2(new_n468), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n473), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n474), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n488), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n500), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n489), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n479), .A2(new_n504), .A3(new_n481), .A4(new_n490), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n492), .A2(new_n503), .A3(new_n286), .A4(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n506), .A2(G472), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n497), .A2(new_n499), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n493), .B1(new_n510), .B2(new_n324), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n511), .B2(new_n501), .ZN(new_n512));
  NOR4_X1   g326(.A1(new_n500), .A2(KEYINPUT31), .A3(new_n493), .A4(new_n488), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n501), .B1(new_n495), .B2(new_n481), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n508), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT30), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n498), .B1(new_n471), .B2(new_n473), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n324), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n475), .A3(new_n501), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT31), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n495), .A2(new_n481), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n488), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n509), .A3(new_n501), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n516), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT71), .B1(new_n507), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n516), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT32), .B1(new_n527), .B2(new_n516), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n506), .A2(G472), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n458), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n485), .A2(new_n277), .A3(G214), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n225), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G131), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(G143), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n258), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(KEYINPUT17), .A3(G131), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n426), .A2(new_n544), .A3(new_n427), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n539), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n417), .A2(new_n421), .A3(new_n422), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n549), .A2(G146), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n431), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n191), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n546), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n540), .A2(new_n542), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(KEYINPUT19), .B2(new_n430), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n427), .B(new_n555), .C1(new_n557), .C2(G146), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n553), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OR3_X1    g376(.A1(new_n560), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT20), .B1(new_n560), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(G234), .A2(G237), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(G952), .A3(new_n277), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(G902), .A3(G953), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT21), .B(G898), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n553), .B1(new_n546), .B2(new_n551), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n286), .B1(new_n554), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G475), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n225), .A2(G128), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n221), .A2(G143), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(KEYINPUT90), .ZN(new_n584));
  INV_X1    g398(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n578), .B2(new_n579), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n250), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G122), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G116), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n316), .A2(G122), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G107), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n189), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n582), .A2(new_n579), .A3(new_n250), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OR3_X1    g413(.A1(new_n590), .A2(KEYINPUT14), .A3(G116), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT91), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n189), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n592), .A2(KEYINPUT14), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n600), .A2(new_n603), .A3(KEYINPUT91), .A4(new_n591), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n250), .B1(new_n582), .B2(new_n579), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n595), .B1(new_n597), .B2(new_n606), .ZN(new_n607));
  OAI22_X1  g421(.A1(new_n589), .A2(new_n599), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n303), .A2(new_n452), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n607), .B1(new_n602), .B2(new_n604), .ZN(new_n613));
  INV_X1    g427(.A(new_n588), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n586), .A2(new_n587), .B1(new_n579), .B2(new_n578), .ZN(new_n615));
  OAI21_X1  g429(.A(G134), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(new_n598), .ZN(new_n617));
  INV_X1    g431(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT93), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n617), .A2(new_n618), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n613), .B(new_n611), .C1(new_n616), .C2(new_n598), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n286), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G478), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(KEYINPUT15), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n621), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n620), .B1(KEYINPUT15), .B2(new_n627), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT94), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n630), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n577), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n407), .A2(new_n537), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT95), .B(G101), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  NAND2_X1  g451(.A1(new_n565), .A2(new_n576), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n618), .B1(new_n608), .B2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n617), .A2(KEYINPUT96), .A3(new_n611), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n622), .B2(new_n623), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n643), .A2(new_n645), .A3(G478), .A4(new_n286), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT97), .B1(new_n639), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n572), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n397), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n404), .A2(new_n405), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT83), .B(new_n305), .C1(new_n401), .C2(new_n403), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n515), .B2(G902), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n527), .A2(new_n516), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n458), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n651), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(new_n633), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n631), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n563), .A2(new_n564), .B1(G475), .B2(new_n575), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n572), .B(KEYINPUT98), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n397), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n654), .A3(new_n658), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NAND2_X1  g483(.A1(new_n429), .A2(new_n435), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n441), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n456), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n449), .B2(new_n454), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n657), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n654), .A2(new_n397), .A3(new_n634), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT37), .B(G110), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G12));
  AOI21_X1  g494(.A(new_n675), .B1(new_n530), .B2(new_n536), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n407), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n569), .A2(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n567), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n686), .A2(new_n662), .A3(new_n631), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(new_n685), .B(KEYINPUT39), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n654), .A2(KEYINPUT40), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT40), .B1(new_n654), .B2(new_n690), .ZN(new_n692));
  OR3_X1    g506(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT102), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT102), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n395), .A2(new_n396), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n632), .A2(new_n638), .A3(new_n307), .A4(new_n633), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n488), .B1(new_n476), .B2(new_n478), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n522), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n286), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n700), .A2(KEYINPUT101), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n533), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n675), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n697), .A2(new_n698), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n693), .A2(new_n694), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  OAI211_X1 g523(.A(new_n638), .B(new_n685), .C1(new_n647), .C2(new_n648), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n683), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  OAI211_X1 g527(.A(new_n401), .B(new_n304), .C1(new_n299), .C2(new_n187), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n651), .A2(new_n537), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND3_X1  g532(.A1(new_n666), .A2(new_n537), .A3(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  AND2_X1   g534(.A1(new_n397), .A2(new_n715), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n681), .A3(new_n634), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AOI21_X1  g537(.A(new_n698), .B1(new_n395), .B2(new_n396), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n523), .A2(new_n526), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n479), .A2(new_n481), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n501), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n479), .A2(KEYINPUT103), .A3(new_n481), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT104), .B1(new_n730), .B2(new_n517), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT69), .B1(new_n493), .B2(new_n494), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n475), .A2(new_n459), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n480), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n481), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n488), .A3(new_n729), .ZN(new_n737));
  INV_X1    g551(.A(new_n725), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n516), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n731), .A2(new_n741), .A3(new_n655), .ZN(new_n742));
  INV_X1    g556(.A(new_n458), .ZN(new_n743));
  INV_X1    g557(.A(new_n665), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n714), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n724), .A2(new_n742), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND4_X1  g561(.A1(new_n731), .A2(new_n741), .A3(new_n655), .A4(new_n674), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n711), .B(new_n721), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NAND2_X1  g566(.A1(new_n528), .A2(KEYINPUT106), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n527), .A2(new_n754), .A3(KEYINPUT32), .A4(new_n516), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n535), .A2(new_n753), .A3(new_n518), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT42), .A3(new_n743), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n404), .A2(new_n307), .A3(new_n395), .A4(new_n396), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n710), .ZN(new_n759));
  INV_X1    g573(.A(new_n758), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n537), .A2(new_n711), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n258), .ZN(G33));
  NAND3_X1  g578(.A1(new_n537), .A2(new_n687), .A3(new_n760), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NOR2_X1   g580(.A1(new_n187), .A2(new_n286), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n402), .A2(KEYINPUT107), .A3(KEYINPUT45), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n285), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n187), .B1(new_n285), .B2(new_n770), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n774), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  INV_X1    g590(.A(new_n401), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n304), .A3(new_n690), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n664), .B1(new_n647), .B2(new_n648), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n664), .C1(new_n647), .C2(new_n648), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n657), .A2(new_n674), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n395), .A2(new_n307), .A3(new_n396), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(new_n787), .A3(new_n785), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n788), .A2(new_n792), .A3(KEYINPUT109), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT109), .B1(new_n788), .B2(new_n792), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n781), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT110), .B(G137), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n304), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n779), .A2(new_n800), .A3(new_n304), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n711), .A2(new_n530), .A3(new_n536), .A4(new_n458), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n789), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NOR3_X1   g619(.A1(new_n458), .A2(new_n308), .A3(new_n305), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT111), .Z(new_n807));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n808));
  INV_X1    g622(.A(new_n299), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n777), .B1(G469), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n705), .A2(new_n782), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n810), .A2(new_n808), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n697), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n801), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n810), .A2(new_n305), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n743), .A2(new_n786), .A3(new_n568), .A4(new_n742), .ZN(new_n819));
  INV_X1    g633(.A(new_n789), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n815), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n821), .B(KEYINPUT116), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n816), .A2(new_n817), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n308), .A3(new_n697), .A4(new_n715), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n749), .A2(new_n750), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n789), .A2(new_n714), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n786), .A2(new_n568), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n705), .A2(new_n458), .A3(new_n567), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n833), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n647), .A2(new_n638), .A3(new_n648), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n832), .A2(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n824), .A2(new_n827), .A3(new_n830), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n743), .A3(new_n756), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n819), .A2(new_n721), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n277), .A2(G952), .ZN(new_n845));
  INV_X1    g659(.A(new_n649), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n825), .A2(new_n826), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n407), .B(new_n681), .C1(new_n687), .C2(new_n711), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n404), .A2(new_n685), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n724), .A2(new_n675), .A3(new_n705), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n751), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n857), .B2(KEYINPUT113), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n306), .A2(new_n397), .A3(new_n406), .A4(new_n634), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n507), .A2(new_n529), .A3(KEYINPUT71), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n743), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n676), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n629), .A2(new_n630), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n649), .B1(new_n873), .B2(new_n638), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n306), .A3(new_n406), .A4(new_n658), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n308), .B(new_n744), .C1(new_n395), .C2(new_n396), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n865), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n654), .A2(new_n658), .A3(new_n876), .A4(new_n874), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n635), .A2(new_n677), .A3(new_n880), .A4(KEYINPUT112), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n716), .A2(new_n719), .A3(new_n722), .A4(new_n746), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n758), .A2(new_n710), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n749), .B2(new_n750), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n686), .A2(new_n872), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n681), .A2(new_n654), .A3(new_n820), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n765), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n763), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n864), .A2(new_n890), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n857), .B(KEYINPUT52), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n882), .A2(new_n889), .A3(new_n883), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n895), .A2(new_n896), .A3(new_n894), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n864), .A2(new_n890), .A3(new_n891), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT115), .B(new_n898), .C1(new_n901), .C2(new_n893), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n898), .A2(KEYINPUT115), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n853), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n814), .B1(new_n904), .B2(new_n905), .ZN(G75));
  XNOR2_X1  g720(.A(new_n356), .B(new_n369), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  NAND2_X1  g722(.A1(G210), .A2(G902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n892), .B2(new_n897), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(KEYINPUT56), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n277), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(KEYINPUT56), .A3(new_n908), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT118), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n910), .A2(KEYINPUT56), .A3(new_n908), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n913), .A4(new_n911), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(new_n767), .B(KEYINPUT57), .ZN(new_n921));
  INV_X1    g735(.A(new_n898), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n893), .B1(new_n892), .B2(new_n897), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n400), .B2(new_n399), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n286), .B1(new_n892), .B2(new_n897), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n772), .A3(new_n773), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n925), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n560), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n912), .ZN(G60));
  NAND2_X1  g747(.A1(new_n643), .A2(new_n645), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n922), .B2(new_n923), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n913), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n902), .A2(new_n903), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n934), .B2(new_n941), .ZN(G63));
  XNOR2_X1  g756(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n452), .A2(new_n286), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n892), .B2(new_n897), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n672), .B(KEYINPUT120), .Z(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n455), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n913), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT61), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n949), .B2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n571), .B2(new_n365), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n882), .A2(new_n883), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(KEYINPUT122), .A3(new_n277), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT122), .B1(new_n959), .B2(new_n277), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n356), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(G898), .B2(new_n277), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT125), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n510), .B(new_n557), .Z(new_n971));
  AND2_X1   g785(.A1(new_n854), .A2(new_n751), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n708), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n820), .A2(new_n874), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n537), .A3(new_n654), .A4(new_n690), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n795), .A2(new_n804), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n708), .A2(new_n978), .A3(new_n972), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n971), .B1(new_n980), .B2(new_n277), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n971), .A2(new_n277), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n724), .A2(new_n743), .A3(new_n756), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n765), .B1(new_n780), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n763), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n795), .A3(new_n804), .A4(new_n972), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n804), .A2(new_n972), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(KEYINPUT123), .A3(new_n795), .A4(new_n985), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n982), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n277), .A2(G900), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n981), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n966), .A2(new_n967), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n970), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n994), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n991), .A2(new_n992), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n996), .B(new_n969), .C1(new_n997), .C2(new_n981), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n980), .B2(new_n959), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n511), .A2(new_n488), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1003), .A2(KEYINPUT127), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT127), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n988), .A2(new_n990), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1002), .B1(new_n1008), .B2(new_n959), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n502), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1004), .ZN(new_n1011));
  INV_X1    g825(.A(new_n502), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n1001), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n901), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1010), .A2(new_n1014), .A3(new_n913), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1007), .A2(new_n1015), .ZN(G57));
endmodule


