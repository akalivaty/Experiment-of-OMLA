//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  AND3_X1   g0026(.A1(new_n215), .A2(new_n225), .A3(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT67), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  AND3_X1   g0047(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT68), .ZN(new_n248));
  AOI21_X1  g0048(.A(KEYINPUT68), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G223), .A3(G1698), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n252), .B(new_n253), .C1(new_n202), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n256), .A3(G274), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n260), .ZN(new_n263));
  INV_X1    g0063(.A(G226), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G169), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(new_n205), .B2(new_n244), .ZN(new_n271));
  NAND4_X1  g0071(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n210), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n211), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n280), .B1(new_n211), .B2(new_n201), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n273), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n271), .A2(new_n210), .A3(new_n285), .A4(new_n272), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n259), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G50), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G50), .B2(new_n285), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n283), .B2(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n258), .A2(new_n293), .A3(new_n266), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n269), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  AOI211_X1 g0097(.A(new_n297), .B(new_n265), .C1(new_n254), .C2(new_n257), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G200), .B2(new_n267), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n284), .B2(new_n291), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n299), .B(new_n305), .C1(new_n300), .C2(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT68), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n246), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n313), .A2(new_n264), .A3(G1698), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n311), .A2(G232), .A3(G1698), .A4(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n257), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n262), .ZN(new_n319));
  INV_X1    g0119(.A(new_n263), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(G238), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G200), .ZN(new_n327));
  INV_X1    g0127(.A(G50), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n278), .A2(new_n328), .B1(new_n211), .B2(G68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n275), .A2(new_n202), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n273), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(new_n285), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT74), .B1(new_n336), .B2(new_n337), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n323), .A2(G190), .A3(new_n325), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n327), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n325), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n324), .B1(new_n318), .B2(new_n321), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n326), .A2(new_n348), .A3(G169), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n349), .C1(new_n293), .C2(new_n326), .ZN(new_n350));
  INV_X1    g0150(.A(new_n341), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n343), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n274), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n288), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n354), .A2(new_n286), .B1(new_n285), .B2(new_n353), .ZN(new_n355));
  AND2_X1   g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n277), .A2(G159), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT75), .B(G20), .C1(new_n356), .C2(new_n357), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT76), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n310), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n244), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n211), .B1(new_n248), .B2(new_n249), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n363), .B1(new_n371), .B2(new_n334), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT3), .B(G33), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT7), .B1(new_n375), .B2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n245), .A2(new_n247), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n370), .A3(new_n211), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(G68), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n363), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n380), .A2(new_n273), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n355), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n264), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n375), .B(new_n383), .C1(G223), .C2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n385), .B(KEYINPUT77), .Z(new_n386));
  AOI21_X1  g0186(.A(new_n256), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G232), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n262), .B1(new_n263), .B2(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n387), .A2(new_n389), .A3(new_n293), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n387), .A2(new_n389), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(G169), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT18), .B1(new_n382), .B2(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n387), .A2(new_n389), .A3(new_n297), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(G200), .B2(new_n391), .ZN(new_n395));
  INV_X1    g0195(.A(new_n355), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n245), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n247), .A3(new_n367), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n311), .B2(new_n312), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT16), .B1(new_n403), .B2(new_n363), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n380), .A2(new_n273), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n395), .B(new_n396), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n396), .B1(new_n404), .B2(new_n405), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  INV_X1    g0210(.A(new_n392), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n374), .A2(new_n381), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n396), .A4(new_n395), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n393), .A2(new_n408), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G244), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n262), .B1(new_n263), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n250), .A2(G238), .A3(G1698), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT72), .B(G107), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n250), .C2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n422), .B2(new_n257), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n293), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n287), .A2(G77), .A3(new_n288), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n275), .B1(new_n211), .B2(new_n202), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n274), .B(KEYINPUT73), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n277), .ZN(new_n430));
  INV_X1    g0230(.A(new_n273), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n426), .B1(G77), .B2(new_n285), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n423), .B2(G169), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(new_n423), .B2(G190), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n423), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n307), .A2(new_n352), .A3(new_n416), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n244), .A2(G1), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n286), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G116), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n285), .A2(G116), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT79), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(G33), .A3(G283), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(G20), .B1(new_n244), .B2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G20), .ZN(new_n454));
  AND4_X1   g0254(.A1(KEYINPUT20), .A2(new_n452), .A3(new_n273), .A4(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n450), .A2(new_n451), .B1(G20), .B2(new_n453), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT20), .B1(new_n456), .B2(new_n273), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n443), .B(new_n445), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(G264), .A2(G1698), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n245), .A2(new_n247), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n375), .A2(new_n462), .A3(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n375), .A2(G257), .A3(new_n251), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n311), .B2(new_n312), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n257), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n256), .ZN(new_n474));
  INV_X1    g0274(.A(G270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n256), .A2(G274), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n468), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n458), .A2(new_n479), .A3(KEYINPUT21), .A4(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(G303), .B1(new_n248), .B2(new_n249), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(new_n463), .A3(new_n464), .A4(new_n461), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(new_n257), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n458), .A2(new_n483), .A3(G179), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n458), .A2(G169), .A3(new_n479), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(G200), .ZN(new_n489));
  INV_X1    g0289(.A(new_n458), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n297), .C2(new_n479), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT72), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G87), .A2(G97), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n211), .B1(new_n316), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n375), .A2(new_n211), .A3(G68), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n275), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(new_n273), .B1(new_n333), .B2(new_n427), .ZN(new_n506));
  INV_X1    g0306(.A(new_n427), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n442), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g0308(.A1(G238), .A2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n417), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n245), .A2(new_n509), .A3(new_n247), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n256), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n256), .A2(G274), .A3(new_n470), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n259), .A2(G45), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n256), .A2(G250), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n506), .A2(new_n508), .B1(new_n293), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n518), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n268), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n273), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n442), .A2(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n427), .A2(new_n333), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n513), .B2(new_n517), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT80), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n506), .A2(KEYINPUT80), .A3(new_n527), .A4(new_n524), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n518), .A2(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n522), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  XOR2_X1   g0333(.A(G97), .B(G107), .Z(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(KEYINPUT6), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n371), .B2(new_n421), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n273), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n285), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n442), .B2(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n542), .A2(new_n417), .A3(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n311), .A2(new_n312), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n311), .A2(G250), .A3(G1698), .A4(new_n312), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n375), .A2(G244), .A3(new_n251), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n542), .B1(new_n449), .B2(new_n447), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n311), .A2(KEYINPUT78), .A3(new_n312), .A4(new_n543), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n257), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n476), .A2(new_n473), .ZN(new_n553));
  INV_X1    g0353(.A(G257), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n474), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n268), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n293), .B(new_n555), .C1(new_n551), .C2(new_n257), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n541), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(G190), .A3(new_n556), .ZN(new_n560));
  INV_X1    g0360(.A(new_n540), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n537), .B2(new_n273), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n551), .B2(new_n257), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n560), .B(new_n562), .C1(new_n437), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n473), .A2(G264), .A3(new_n256), .ZN(new_n565));
  XOR2_X1   g0365(.A(KEYINPUT83), .B(G294), .Z(new_n566));
  NOR2_X1   g0366(.A1(new_n251), .A2(G257), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G250), .A2(G1698), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(G33), .A2(new_n566), .B1(new_n569), .B2(new_n375), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n553), .B(new_n565), .C1(new_n570), .C2(new_n256), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n268), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n377), .A2(new_n568), .A3(new_n567), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT83), .B(G294), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n244), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n257), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n293), .A3(new_n553), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n421), .B2(G20), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n493), .A3(G20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n453), .C2(new_n275), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G87), .ZN(new_n586));
  OR3_X1    g0386(.A1(new_n586), .A2(KEYINPUT22), .A3(G20), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n248), .A2(new_n249), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n245), .A2(new_n247), .A3(new_n211), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n585), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n313), .B2(new_n587), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n593), .A3(new_n585), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n431), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n442), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n493), .ZN(new_n600));
  INV_X1    g0400(.A(G13), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(G1), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G20), .A3(new_n493), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT25), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n579), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n592), .A2(new_n594), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n593), .B1(new_n596), .B2(new_n585), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n273), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n576), .A2(new_n297), .A3(new_n553), .A4(new_n565), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n611), .A2(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n571), .A2(new_n437), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(KEYINPUT84), .A3(new_n611), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n610), .A2(new_n605), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n559), .A2(new_n564), .A3(new_n607), .A4(new_n615), .ZN(new_n616));
  NOR4_X1   g0416(.A1(new_n440), .A2(new_n492), .A3(new_n532), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n343), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n434), .B1(new_n350), .B2(new_n351), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n408), .A2(new_n414), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n393), .B(new_n412), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n304), .A2(new_n306), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n296), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n440), .ZN(new_n624));
  INV_X1    g0424(.A(new_n513), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT85), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT85), .B1(new_n514), .B2(new_n516), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n268), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n519), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT26), .B1(new_n559), .B2(new_n532), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT86), .B1(new_n557), .B2(new_n558), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n552), .A2(G179), .A3(new_n556), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT86), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n633), .B(new_n634), .C1(new_n268), .C2(new_n563), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n530), .A2(new_n506), .A3(new_n524), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n628), .A2(G200), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n519), .B2(new_n629), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n632), .A2(new_n635), .A3(new_n541), .A4(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n630), .B(new_n631), .C1(new_n639), .C2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT87), .ZN(new_n641));
  INV_X1    g0441(.A(new_n630), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n633), .B1(new_n268), .B2(new_n563), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT80), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n506), .A2(new_n524), .ZN(new_n645));
  INV_X1    g0445(.A(new_n527), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n530), .A3(new_n529), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n643), .A2(new_n648), .A3(new_n522), .A4(new_n541), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(KEYINPUT26), .C2(new_n639), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n559), .A2(new_n564), .A3(new_n615), .A4(new_n638), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n578), .B1(new_n610), .B2(new_n605), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n483), .A2(new_n268), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT21), .B1(new_n655), .B2(new_n458), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n480), .A2(new_n484), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n641), .A2(new_n652), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n624), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n623), .A2(new_n662), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n485), .A2(new_n488), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n602), .A2(new_n211), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(KEYINPUT88), .A3(KEYINPUT27), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT88), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(G213), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n490), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n676), .B(KEYINPUT89), .C1(new_n492), .C2(new_n675), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n664), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n615), .A2(new_n607), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n673), .B1(new_n598), .B2(new_n606), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n654), .A2(new_n673), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n607), .A2(new_n673), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n673), .B1(new_n485), .B2(new_n488), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n683), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n498), .A2(G116), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n206), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n694), .A2(new_n259), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n214), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NAND2_X1  g0499(.A1(new_n661), .A2(new_n674), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n659), .B1(new_n640), .B2(KEYINPUT87), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n673), .B1(new_n704), .B2(new_n652), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT91), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n630), .B1(new_n649), .B2(KEYINPUT26), .C1(new_n653), .C2(new_n658), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT29), .B(new_n674), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n468), .A2(G179), .A3(new_n478), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n518), .A2(new_n565), .A3(new_n576), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n563), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n563), .A2(new_n711), .A3(KEYINPUT30), .A4(new_n712), .ZN(new_n716));
  INV_X1    g0516(.A(new_n563), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n628), .A2(new_n571), .A3(new_n293), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n479), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n673), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR4_X1   g0525(.A1(new_n616), .A2(new_n492), .A3(new_n532), .A4(new_n673), .ZN(new_n726));
  OAI21_X1  g0526(.A(G330), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n720), .B2(new_n673), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n616), .ZN(new_n732));
  INV_X1    g0532(.A(new_n492), .ZN(new_n733));
  INV_X1    g0533(.A(new_n532), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .A4(new_n674), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT90), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n728), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n710), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n601), .A2(G20), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n259), .A3(new_n696), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n682), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n677), .A2(new_n679), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n745), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n297), .A2(new_n437), .ZN(new_n757));
  NAND2_X1  g0557(.A1(G20), .A2(G179), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(G190), .A3(new_n437), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n211), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n762), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G322), .A2(new_n767), .B1(new_n770), .B2(G329), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n437), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n759), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI221_X1 g0576(.A(new_n771), .B1(new_n772), .B2(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n211), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n765), .B(new_n777), .C1(new_n566), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n757), .A2(new_n768), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n313), .B1(new_n466), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  INV_X1    g0584(.A(new_n782), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G87), .A2(new_n785), .B1(new_n767), .B2(G58), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n780), .A2(G97), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n786), .A2(new_n250), .A3(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n774), .A2(new_n493), .B1(new_n763), .B2(new_n202), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n760), .A2(new_n328), .B1(new_n775), .B2(new_n334), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n769), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n770), .A2(KEYINPUT32), .A3(G159), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n789), .B(new_n790), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n781), .A2(new_n784), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n210), .B1(G20), .B2(new_n268), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n752), .A2(new_n797), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n250), .A2(G355), .A3(new_n206), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n242), .A2(new_n469), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n695), .A2(new_n375), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n213), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n801), .B1(G116), .B2(new_n206), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n756), .B(new_n799), .C1(new_n800), .C2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n746), .A2(new_n749), .B1(new_n755), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  INV_X1    g0608(.A(KEYINPUT95), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n425), .B2(new_n433), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n422), .A2(new_n257), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n268), .B1(new_n811), .B2(new_n418), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n812), .A2(KEYINPUT95), .A3(new_n424), .A4(new_n432), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n673), .A2(new_n432), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n813), .A3(new_n438), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n434), .A2(new_n673), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n700), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n810), .A2(new_n813), .A3(new_n438), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n661), .A2(new_n674), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n739), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n818), .A2(new_n728), .A3(new_n738), .A4(new_n820), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n823), .A3(new_n756), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n797), .A2(new_n750), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n745), .B1(G77), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n782), .A2(new_n493), .B1(new_n769), .B2(new_n764), .ZN(new_n828));
  INV_X1    g0628(.A(new_n760), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G303), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n766), .A2(new_n831), .B1(new_n774), .B2(new_n586), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n775), .A2(new_n772), .B1(new_n763), .B2(new_n453), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n830), .A2(new_n313), .A3(new_n787), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n760), .A2(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n775), .A2(new_n276), .B1(new_n763), .B2(new_n792), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(G143), .C2(new_n767), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n377), .B1(new_n770), .B2(G132), .ZN(new_n841));
  INV_X1    g0641(.A(G58), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n779), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n774), .A2(new_n334), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G50), .B2(new_n785), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT94), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT34), .B2(new_n839), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n835), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n827), .B1(new_n848), .B2(new_n797), .ZN(new_n849));
  INV_X1    g0649(.A(new_n817), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n751), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n824), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT97), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT97), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n824), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(G384));
  OR2_X1    g0657(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(G116), .A3(new_n212), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n214), .B(G77), .C1(new_n842), .C2(new_n334), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n328), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n259), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n409), .A2(new_n411), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n409), .A2(new_n670), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(new_n406), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n866), .A2(new_n867), .A3(new_n870), .A4(new_n406), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n415), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT98), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n363), .A2(new_n379), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n381), .B1(KEYINPUT16), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n671), .B1(new_n881), .B2(new_n396), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n415), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n406), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n881), .A2(new_n396), .B1(new_n392), .B2(new_n671), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n871), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n869), .A2(new_n871), .B1(new_n415), .B2(new_n873), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n888), .B(new_n879), .C1(new_n890), .C2(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT98), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n883), .A2(new_n887), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n876), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n879), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n350), .A2(new_n351), .A3(new_n674), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n346), .A2(KEYINPUT14), .B1(new_n326), .B2(new_n293), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n348), .B1(new_n326), .B2(G169), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n351), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n351), .A2(new_n673), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n618), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n351), .B(new_n673), .C1(new_n350), .C2(new_n343), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n810), .A2(new_n813), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n674), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n820), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n894), .A2(new_n888), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n393), .A2(new_n412), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n671), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n898), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n703), .A2(new_n706), .A3(new_n624), .A4(new_n709), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n623), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n877), .A2(new_n888), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n817), .B1(new_n903), .B2(new_n904), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n736), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT40), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n919), .A2(new_n736), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT40), .B1(new_n894), .B2(new_n888), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n440), .B1(new_n735), .B2(new_n731), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n681), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n925), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n259), .B2(new_n742), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n917), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n865), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NAND4_X1  g0732(.A1(new_n632), .A2(new_n635), .A3(new_n541), .A4(new_n673), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n541), .A2(new_n673), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n559), .A2(new_n564), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n674), .B1(new_n656), .B2(new_n657), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n615), .A2(new_n607), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n933), .A2(new_n935), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n559), .B1(new_n943), .B2(new_n607), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n674), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n674), .A2(new_n526), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n630), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n638), .B2(new_n947), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT99), .Z(new_n950));
  XNOR2_X1  g0750(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n946), .B(new_n952), .C1(new_n953), .C2(new_n950), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n946), .B2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(new_n687), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n680), .A2(new_n681), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n936), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n955), .B(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n744), .A2(new_n259), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT45), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT101), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n691), .A2(new_n963), .A3(new_n936), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(new_n691), .B2(new_n936), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n937), .A2(new_n938), .B1(new_n607), .B2(new_n673), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT101), .B1(new_n943), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n691), .A2(new_n963), .A3(new_n936), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n943), .A2(KEYINPUT44), .A3(new_n967), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n691), .B2(new_n936), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n966), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n957), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n688), .A2(new_n966), .A3(new_n970), .A4(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n956), .A2(new_n937), .ZN(new_n979));
  INV_X1    g0779(.A(new_n939), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT102), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n747), .B2(G330), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n681), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n980), .B(new_n979), .C1(new_n682), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n739), .B(new_n710), .C1(new_n978), .C2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n696), .B(KEYINPUT41), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT103), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n961), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(KEYINPUT103), .A3(new_n989), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n959), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n950), .A2(new_n752), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n800), .B1(new_n206), .B2(new_n427), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n235), .B2(new_n803), .ZN(new_n997));
  INV_X1    g0797(.A(new_n775), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n566), .A2(new_n998), .B1(new_n770), .B2(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n764), .B2(new_n760), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n782), .B2(new_n453), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(new_n421), .C2(new_n779), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n377), .B1(new_n763), .B2(new_n772), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n766), .A2(new_n466), .B1(new_n774), .B2(new_n503), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1000), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n763), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n767), .A2(G150), .B1(new_n1008), .B2(G50), .ZN(new_n1009));
  INV_X1    g0809(.A(G143), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n760), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n780), .A2(G68), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n250), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n774), .A2(new_n202), .B1(new_n769), .B2(new_n836), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n782), .A2(new_n842), .B1(new_n775), .B2(new_n792), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  AOI211_X1 g0818(.A(new_n756), .B(new_n997), .C1(new_n1018), .C2(new_n797), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n995), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n994), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(G317), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n766), .A2(new_n1024), .B1(new_n763), .B2(new_n466), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT104), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(KEYINPUT104), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G322), .A2(new_n829), .B1(new_n998), .B2(G311), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT105), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n780), .A2(G283), .B1(new_n785), .B2(new_n566), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n377), .B1(new_n769), .B2(new_n761), .C1(new_n453), .C2(new_n774), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n760), .A2(new_n792), .B1(new_n775), .B2(new_n274), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n774), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n377), .B(new_n1041), .C1(G97), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n780), .A2(new_n507), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n769), .A2(new_n276), .B1(new_n763), .B2(new_n334), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n202), .A2(new_n782), .B1(new_n766), .B2(new_n328), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n797), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n694), .A2(new_n206), .A3(new_n250), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n232), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n803), .B1(new_n1051), .B2(new_n469), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n429), .A2(new_n328), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n469), .B1(new_n334), .B2(new_n202), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n694), .A3(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1050), .B1(G107), .B2(new_n206), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n756), .B1(new_n1057), .B2(new_n800), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1049), .B(new_n1058), .C1(new_n687), .C2(new_n753), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT106), .Z(new_n1060));
  INV_X1    g0860(.A(new_n987), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n739), .A3(new_n710), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n696), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n740), .A2(new_n1061), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1060), .B1(new_n987), .B2(new_n960), .C1(new_n1063), .C2(new_n1064), .ZN(G393));
  INV_X1    g0865(.A(new_n978), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n961), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n800), .B1(new_n503), .B2(new_n206), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n239), .B2(new_n803), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G283), .A2(new_n785), .B1(new_n770), .B2(G322), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT107), .Z(new_n1071));
  OAI22_X1  g0871(.A1(new_n774), .A2(new_n493), .B1(new_n763), .B2(new_n831), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G303), .B2(new_n998), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n250), .B1(G116), .B2(new_n780), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1024), .A2(new_n760), .B1(new_n766), .B2(new_n764), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n276), .A2(new_n760), .B1(new_n766), .B2(new_n792), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n782), .A2(new_n334), .B1(new_n769), .B2(new_n1010), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G50), .B2(new_n998), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n429), .A2(new_n1008), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n779), .A2(new_n202), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n377), .B1(new_n1042), .B2(G87), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1075), .A2(new_n1077), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n756), .B(new_n1069), .C1(new_n1087), .C2(new_n797), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n936), .B2(new_n753), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1061), .A2(new_n739), .A3(new_n710), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(new_n1066), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n696), .B1(new_n1062), .B2(new_n978), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1067), .B(new_n1089), .C1(new_n1091), .C2(new_n1092), .ZN(G390));
  INV_X1    g0893(.A(new_n696), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n897), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n896), .B1(new_n909), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n674), .B(new_n819), .C1(new_n707), .C2(new_n708), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n908), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n897), .B(new_n918), .C1(new_n1099), .C2(new_n906), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n728), .A2(new_n738), .A3(new_n919), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1096), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n918), .A2(new_n897), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n905), .B2(new_n1098), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n705), .A2(new_n819), .B1(new_n674), .B2(new_n907), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n897), .B1(new_n1105), .B2(new_n906), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n896), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n681), .B1(new_n731), .B2(new_n735), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n919), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1102), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n624), .A2(new_n1108), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n915), .A2(new_n623), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n728), .A2(new_n738), .A3(new_n850), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1113), .A2(new_n906), .B1(new_n1108), .B2(new_n919), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n817), .B1(new_n727), .B2(KEYINPUT108), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT108), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n905), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1114), .A2(new_n1105), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1094), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT109), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1096), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1109), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1113), .A2(new_n906), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1109), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1105), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n906), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n915), .A2(new_n623), .A3(new_n1111), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1110), .A2(new_n1121), .A3(KEYINPUT109), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1122), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n896), .A2(new_n750), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n745), .B1(new_n353), .B2(new_n826), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n782), .A2(new_n586), .B1(new_n774), .B2(new_n334), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n760), .A2(new_n772), .B1(new_n763), .B2(new_n503), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n250), .A2(new_n1141), .A3(new_n1083), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n421), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G116), .A2(new_n767), .B1(new_n998), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n831), .C2(new_n769), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT111), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n760), .A2(new_n1149), .B1(new_n763), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n785), .A2(G150), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1152), .A2(KEYINPUT53), .B1(new_n792), .B2(new_n779), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(KEYINPUT53), .C2(new_n1152), .ZN(new_n1154));
  INV_X1    g0954(.A(G132), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n766), .A2(new_n1155), .B1(new_n769), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n998), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n313), .B1(G50), .B2(new_n1042), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT110), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1148), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1140), .B1(new_n1163), .B2(new_n797), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1126), .A2(new_n961), .B1(new_n1139), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1138), .A2(new_n1165), .ZN(G378));
  AOI22_X1  g0966(.A1(new_n829), .A2(G116), .B1(new_n770), .B2(G283), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n842), .B2(new_n774), .C1(new_n493), .C2(new_n766), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n427), .A2(new_n763), .B1(new_n775), .B2(new_n503), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT112), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n375), .A2(G41), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1012), .B(new_n1171), .C1(new_n202), .C2(new_n782), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT113), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(G33), .A2(G41), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1171), .A2(G50), .A3(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1156), .A2(new_n760), .B1(new_n766), .B2(new_n1149), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G137), .B2(new_n1008), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1150), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n785), .A2(new_n1180), .B1(new_n998), .B2(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n276), .C2(new_n779), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  INV_X1    g0983(.A(G124), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1176), .B1(new_n769), .B2(new_n1184), .C1(new_n792), .C2(new_n774), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1182), .B2(KEYINPUT59), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1175), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n797), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT114), .Z(new_n1191));
  AOI211_X1 g0991(.A(new_n756), .B(new_n1191), .C1(new_n328), .C2(new_n825), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n292), .A2(new_n670), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n307), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n307), .A2(new_n1193), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n750), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1192), .A2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n920), .A2(KEYINPUT40), .B1(new_n922), .B2(new_n923), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1202), .B1(new_n1205), .B2(new_n681), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n925), .A2(G330), .A3(new_n1201), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(KEYINPUT115), .A3(new_n914), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n914), .B1(new_n1208), .B2(KEYINPUT115), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1212), .B2(new_n960), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1112), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1211), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1209), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1208), .B(new_n914), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT57), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1126), .A2(new_n1123), .A3(new_n1135), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT109), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1134), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n696), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1214), .B1(new_n1218), .B2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1121), .A3(new_n989), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT116), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n960), .B(KEYINPUT117), .Z(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n906), .A2(new_n750), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n745), .B1(G68), .B2(new_n826), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n831), .A2(new_n760), .B1(new_n766), .B2(new_n772), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1144), .B2(new_n1008), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n782), .A2(new_n503), .B1(new_n775), .B2(new_n453), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n774), .A2(new_n202), .B1(new_n769), .B2(new_n466), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n313), .A3(new_n1044), .A4(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n769), .A2(new_n1149), .B1(new_n763), .B2(new_n276), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n375), .B1(new_n774), .B2(new_n842), .C1(new_n779), .C2(new_n328), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(G159), .C2(new_n785), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT118), .Z(new_n1242));
  AOI22_X1  g1042(.A1(G137), .A2(new_n767), .B1(new_n998), .B2(new_n1180), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1155), .B2(new_n760), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1238), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1232), .B1(new_n1245), .B2(new_n797), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1120), .A2(new_n1230), .B1(new_n1231), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1228), .A2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT57), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1208), .A2(new_n914), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1208), .A2(new_n914), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1094), .B1(new_n1215), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1252), .B1(new_n1223), .B2(new_n1212), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1213), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G381), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1251), .A2(new_n1258), .A3(new_n1022), .A4(new_n1259), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n672), .A2(G213), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT119), .Z(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1249), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G407), .A2(G213), .A3(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G393), .B(new_n807), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n994), .B2(new_n1021), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n988), .A2(KEYINPUT103), .A3(new_n989), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT103), .B1(new_n988), .B2(new_n989), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n961), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1020), .B(G390), .C1(new_n1271), .C2(new_n959), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT124), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1277), .A3(new_n1274), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1266), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1280));
  AOI211_X1 g1080(.A(KEYINPUT124), .B(KEYINPUT125), .C1(new_n1268), .C2(new_n1272), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1266), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1265), .B1(new_n1279), .B2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1214), .C1(new_n1218), .C2(new_n1224), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1215), .A2(new_n989), .A3(new_n1217), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1219), .A2(new_n1230), .B1(new_n1203), .B2(new_n1192), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1249), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1262), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1094), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT120), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1133), .A2(new_n1295), .A3(KEYINPUT60), .A4(new_n1134), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1134), .A3(KEYINPUT60), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT120), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1294), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1247), .ZN(new_n1302));
  OAI21_X1  g1102(.A(G384), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1296), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n696), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT60), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G384), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1247), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT63), .B1(new_n1290), .B2(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1284), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1262), .A2(G2897), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1309), .B1(new_n1308), .B2(new_n1247), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1302), .B(G384), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT121), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT121), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1311), .A2(new_n1319), .A3(new_n1314), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1314), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1303), .A2(new_n1310), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT122), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1303), .A2(KEYINPUT122), .A3(new_n1310), .A4(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1321), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT123), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1290), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT123), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1321), .A2(new_n1327), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(G378), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1334), .B1(new_n1258), .B2(G378), .ZN(new_n1335));
  OAI21_X1  g1135(.A(KEYINPUT126), .B1(new_n1335), .B2(new_n1262), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1262), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1336), .A2(new_n1340), .A3(KEYINPUT63), .A4(new_n1311), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1313), .A2(new_n1333), .A3(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(new_n1336), .A2(new_n1340), .B1(new_n1328), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1290), .A2(new_n1344), .A3(new_n1311), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1311), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT61), .B1(new_n1347), .B2(KEYINPUT62), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1343), .B1(new_n1345), .B2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1342), .A2(new_n1350), .ZN(G405));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1249), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1353), .A2(new_n1285), .A3(new_n1347), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1347), .B1(new_n1353), .B2(new_n1285), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1352), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1285), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1311), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1353), .A2(new_n1285), .A3(new_n1347), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(KEYINPUT127), .A3(new_n1359), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1356), .B(new_n1360), .C1(new_n1283), .C2(new_n1279), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1343), .B(new_n1352), .C1(new_n1355), .C2(new_n1354), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


