//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G110), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n194), .B(KEYINPUT72), .Z(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  OR2_X1    g011(.A1(G125), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(G125), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n201), .B(G146), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n203), .A2(new_n204), .B1(G119), .B2(new_n191), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(new_n202), .A3(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n205), .A2(new_n206), .B1(new_n193), .B2(G110), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT22), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT73), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n213), .A3(new_n219), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(G234), .B2(new_n224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(G902), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT74), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT32), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT31), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n188), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n218), .A2(KEYINPUT11), .A3(G134), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n249), .A2(new_n250), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n218), .A2(G134), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n248), .A2(G137), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n211), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n259), .B(G146), .C1(new_n191), .C2(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n191), .A2(new_n211), .A3(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n253), .B(new_n256), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n249), .A2(new_n252), .A3(new_n250), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n253), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n260), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n258), .A2(new_n260), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n246), .A2(new_n265), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n262), .A3(new_n263), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT65), .A3(new_n253), .A4(new_n256), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n245), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n265), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n275), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n278), .A2(KEYINPUT64), .A3(new_n253), .A4(new_n256), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n245), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n244), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n265), .A2(new_n246), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n283), .A3(new_n279), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n244), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(G101), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT66), .A2(G237), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT66), .A2(G237), .ZN(new_n294));
  AOI21_X1  g108(.A(G953), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G210), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n292), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n288), .A2(KEYINPUT30), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n282), .A2(new_n283), .A3(new_n245), .A4(new_n284), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n289), .B1(new_n302), .B2(new_n244), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n297), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n237), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n286), .A2(new_n237), .A3(new_n290), .A4(new_n297), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n303), .A2(new_n309), .A3(new_n237), .A4(new_n297), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n244), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT28), .B1(new_n313), .B2(new_n289), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n283), .A2(new_n243), .A3(new_n265), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n313), .C2(new_n289), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n297), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n306), .A2(new_n311), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G472), .A2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n236), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n304), .B1(new_n303), .B2(new_n297), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n304), .A2(new_n286), .A3(new_n290), .A4(new_n297), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT31), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n320), .ZN(new_n329));
  INV_X1    g143(.A(new_n297), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n328), .A2(new_n331), .A3(new_n308), .A4(new_n310), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT32), .A3(new_n323), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(KEYINPUT70), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n335), .A3(KEYINPUT32), .A4(new_n323), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G472), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n303), .A2(new_n297), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(new_n340), .C1(new_n329), .C2(new_n330), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n288), .B(new_n244), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n318), .B1(new_n342), .B2(KEYINPUT28), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n330), .A2(new_n339), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n338), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n235), .B1(new_n337), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G475), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n295), .A2(G143), .A3(G214), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT66), .A2(G237), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT66), .A2(G237), .ZN(new_n354));
  OAI211_X1 g168(.A(G214), .B(new_n215), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n259), .ZN(new_n356));
  AOI211_X1 g170(.A(new_n351), .B(new_n251), .C1(new_n352), .C2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n350), .B1(new_n357), .B2(new_n202), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n201), .B(new_n211), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n251), .B1(new_n352), .B2(new_n356), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n359), .B(KEYINPUT88), .C1(new_n361), .C2(new_n351), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n352), .A2(new_n251), .A3(new_n356), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n351), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n358), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(G104), .Z(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT18), .A2(G131), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(new_n356), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n200), .A2(KEYINPUT85), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n198), .A2(new_n371), .A3(new_n199), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT86), .B(new_n211), .C1(new_n370), .C2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n212), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n372), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(G146), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n376), .B2(KEYINPUT86), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n360), .A2(KEYINPUT84), .A3(KEYINPUT18), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n360), .B2(KEYINPUT18), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n369), .B(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n365), .A2(new_n367), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n363), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n200), .ZN(new_n384));
  INV_X1    g198(.A(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI221_X1 g201(.A(new_n210), .B1(new_n382), .B2(new_n360), .C1(new_n387), .C2(G146), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n367), .B1(new_n380), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n349), .B(new_n224), .C1(new_n381), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT20), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n380), .A2(new_n388), .ZN(new_n392));
  INV_X1    g206(.A(new_n367), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n365), .A2(new_n367), .A3(new_n380), .ZN(new_n395));
  AOI21_X1  g209(.A(G475), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n224), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G217), .A3(new_n215), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n405), .A2(KEYINPUT91), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(KEYINPUT91), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G128), .B(G143), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n248), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n410), .A2(new_n412), .B1(new_n248), .B2(new_n409), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT90), .B(G122), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  INV_X1    g229(.A(G122), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G116), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G107), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n415), .B2(new_n418), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n413), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n424), .A3(G107), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n409), .B(new_n248), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n415), .B(new_n418), .C1(KEYINPUT14), .C2(new_n421), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n408), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n406), .A2(new_n428), .A3(new_n423), .A4(new_n407), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n224), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n401), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(KEYINPUT92), .A3(new_n224), .A4(new_n431), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n434), .B1(new_n437), .B2(new_n401), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G952), .A3(new_n215), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G898), .Z(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n367), .B1(new_n365), .B2(new_n380), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n224), .B1(new_n381), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT89), .B(G475), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n399), .A2(new_n438), .A3(new_n443), .A4(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n404), .A2(new_n224), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(G221), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT3), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n421), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT3), .A2(G107), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(G104), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G101), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT76), .B(G104), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(G104), .A2(G107), .ZN(new_n460));
  OAI211_X1 g274(.A(G101), .B(new_n460), .C1(new_n458), .C2(G107), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n278), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT10), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n458), .A2(new_n455), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n455), .A2(G104), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n453), .B2(new_n421), .ZN(new_n468));
  OAI21_X1  g282(.A(G101), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n469), .A3(KEYINPUT4), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(G101), .C1(new_n466), .C2(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n275), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT10), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n462), .B2(new_n463), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n268), .ZN(new_n477));
  INV_X1    g291(.A(new_n268), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n465), .A2(new_n473), .A3(new_n478), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G140), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n215), .A2(G227), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n481), .B(new_n482), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT79), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n278), .B1(new_n459), .B2(new_n461), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n464), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT77), .B(KEYINPUT12), .C1(new_n488), .C2(new_n478), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n462), .B(new_n463), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n491));
  OR2_X1    g305(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n268), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n489), .A2(new_n493), .A3(new_n483), .A4(new_n479), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n486), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(new_n486), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n224), .ZN(new_n498));
  AND4_X1   g312(.A1(new_n484), .A2(new_n489), .A3(new_n493), .A4(new_n479), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n484), .B1(new_n477), .B2(new_n479), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT78), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n480), .A2(new_n483), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n489), .A2(new_n493), .A3(new_n484), .A4(new_n479), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n505), .A3(G469), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n497), .A2(new_n224), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G214), .B1(G237), .B2(G902), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT80), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n275), .A2(G125), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(G125), .B2(new_n463), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n215), .A2(G224), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n518));
  INV_X1    g332(.A(new_n238), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(G113), .C1(new_n241), .C2(new_n518), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n241), .A2(new_n242), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n462), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n470), .A2(new_n244), .A3(new_n472), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G110), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n528), .A3(new_n526), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n517), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT6), .B1(new_n527), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n516), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n514), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n523), .A2(new_n462), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n520), .A2(G113), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n524), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n528), .B(KEYINPUT8), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n531), .B(new_n536), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n534), .A2(new_n224), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n534), .A2(new_n224), .A3(new_n547), .A4(new_n549), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n512), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n449), .A2(new_n452), .A3(new_n509), .A4(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n348), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G101), .ZN(G3));
  OAI21_X1  g371(.A(G472), .B1(new_n322), .B2(G902), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n324), .B2(new_n322), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n509), .A2(new_n452), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n559), .A2(new_n560), .A3(new_n235), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n391), .A2(new_n398), .B1(new_n445), .B2(new_n446), .ZN(new_n562));
  INV_X1    g376(.A(new_n432), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G478), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n430), .A2(new_n431), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n429), .A2(KEYINPUT93), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT33), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n430), .A2(new_n566), .A3(KEYINPUT33), .A4(new_n431), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n564), .B1(new_n570), .B2(G478), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n510), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n551), .B2(new_n552), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n443), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n561), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT34), .B(G104), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G6));
  XNOR2_X1  g392(.A(new_n447), .B(KEYINPUT94), .ZN(new_n579));
  INV_X1    g393(.A(new_n438), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n399), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n551), .A2(new_n552), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n510), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n443), .B(KEYINPUT95), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n561), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G107), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G9));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n220), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(new_n214), .Z(new_n591));
  AOI22_X1  g405(.A1(new_n227), .A2(new_n229), .B1(new_n233), .B2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n554), .A2(new_n559), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT37), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G110), .ZN(G12));
  NAND2_X1  g409(.A1(new_n337), .A2(new_n347), .ZN(new_n596));
  INV_X1    g410(.A(new_n592), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n440), .B1(new_n442), .B2(G900), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n509), .A2(new_n452), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n599), .A2(new_n581), .A3(new_n583), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G128), .ZN(G30));
  NAND2_X1  g416(.A1(new_n399), .A2(new_n447), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n598), .B(KEYINPUT39), .Z(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n509), .A2(new_n452), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n580), .B(new_n603), .C1(new_n606), .C2(KEYINPUT40), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n551), .A2(new_n552), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT38), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n299), .A2(new_n305), .B1(new_n330), .B2(new_n342), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n611), .B2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n337), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n573), .B1(new_n606), .B2(KEYINPUT40), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n610), .A2(new_n592), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G143), .ZN(G45));
  NOR2_X1   g430(.A1(new_n599), .A2(new_n583), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n596), .A2(new_n572), .A3(new_n597), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G146), .ZN(G48));
  NAND2_X1  g433(.A1(new_n495), .A2(new_n496), .ZN(new_n620));
  OAI21_X1  g434(.A(G469), .B1(new_n620), .B2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n452), .A3(new_n498), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n348), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n575), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT41), .B(G113), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G15));
  NAND3_X1  g442(.A1(new_n348), .A2(new_n585), .A3(new_n623), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n348), .A2(KEYINPUT97), .A3(new_n585), .A4(new_n623), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G116), .ZN(G18));
  AOI21_X1  g448(.A(new_n592), .B1(new_n337), .B2(new_n347), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n622), .A2(new_n583), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n449), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G119), .ZN(G21));
  AOI21_X1  g452(.A(new_n338), .B1(new_n332), .B2(new_n224), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n323), .B(KEYINPUT98), .Z(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n306), .A2(new_n311), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n343), .A2(new_n297), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n235), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n603), .A2(new_n580), .A3(KEYINPUT99), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n562), .B2(new_n438), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n650), .A3(new_n574), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n647), .A2(new_n651), .A3(new_n584), .A4(new_n622), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n416), .ZN(G24));
  INV_X1    g467(.A(new_n598), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n562), .A2(new_n571), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n642), .A2(new_n643), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n640), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n655), .A2(new_n597), .A3(new_n558), .A4(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n574), .A2(new_n452), .A3(new_n498), .A4(new_n621), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT100), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n639), .A2(new_n592), .A3(new_n644), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n636), .A2(new_n661), .A3(new_n662), .A4(new_n655), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G125), .ZN(G27));
  OAI21_X1  g479(.A(G469), .B1(new_n499), .B2(new_n500), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT101), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n668), .B(G469), .C1(new_n499), .C2(new_n500), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n498), .A2(new_n667), .A3(new_n508), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .A3(new_n452), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT102), .B1(new_n670), .B2(new_n452), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n608), .A2(new_n510), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n325), .A2(new_n347), .A3(new_n333), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n646), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n655), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT42), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n348), .A2(new_n681), .A3(new_n675), .A4(new_n598), .ZN(new_n682));
  INV_X1    g496(.A(new_n572), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n251), .ZN(G33));
  INV_X1    g499(.A(new_n581), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n348), .A2(new_n686), .A3(new_n675), .A4(new_n598), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT103), .B(G134), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G36));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n501), .B2(new_n505), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n693), .A2(new_n694), .A3(new_n497), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT45), .B1(new_n499), .B2(new_n500), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n694), .B1(new_n693), .B2(new_n497), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n696), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n691), .B(new_n692), .C1(new_n703), .C2(new_n507), .ZN(new_n704));
  INV_X1    g518(.A(new_n498), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n507), .B1(new_n700), .B2(new_n701), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT106), .B1(new_n706), .B2(KEYINPUT46), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n452), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n690), .B1(new_n710), .B2(new_n604), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n562), .B(KEYINPUT108), .ZN(new_n712));
  INV_X1    g526(.A(new_n571), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT43), .ZN(new_n715));
  OR3_X1    g529(.A1(new_n603), .A2(KEYINPUT43), .A3(new_n571), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n559), .A2(new_n715), .A3(new_n597), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT109), .B1(new_n717), .B2(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n674), .B1(new_n717), .B2(KEYINPUT44), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n452), .A4(new_n605), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n711), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G137), .ZN(G39));
  NOR3_X1   g542(.A1(new_n596), .A2(new_n683), .A3(new_n654), .ZN(new_n729));
  INV_X1    g543(.A(new_n674), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n235), .A3(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(KEYINPUT110), .Z(new_n732));
  NAND3_X1  g546(.A1(new_n709), .A2(KEYINPUT47), .A3(new_n452), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT47), .B1(new_n709), .B2(new_n452), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT111), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G140), .ZN(G42));
  NAND2_X1  g552(.A1(new_n621), .A2(new_n498), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT112), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT49), .Z(new_n741));
  NOR4_X1   g555(.A1(new_n741), .A2(new_n451), .A3(new_n512), .A4(new_n714), .ZN(new_n742));
  INV_X1    g556(.A(new_n613), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n646), .A3(new_n743), .A4(new_n609), .ZN(new_n744));
  INV_X1    g558(.A(new_n735), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n451), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n733), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n440), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n715), .A2(new_n748), .A3(new_n716), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n647), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n747), .A2(new_n730), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n674), .A2(new_n622), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(new_n661), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n743), .A2(new_n646), .A3(new_n748), .A4(new_n755), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n562), .A3(new_n571), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT118), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n609), .A2(new_n573), .A3(new_n623), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT117), .Z(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n752), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT50), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n754), .A2(new_n756), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n637), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n631), .B2(new_n632), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n652), .B1(new_n624), .B2(new_n575), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n670), .A2(new_n452), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n651), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n613), .A2(new_n592), .A3(new_n598), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n618), .A2(new_n778), .A3(new_n601), .A4(new_n664), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n635), .A2(new_n600), .B1(new_n660), .B2(new_n663), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT52), .A3(new_n618), .A4(new_n778), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n781), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT115), .B1(new_n781), .B2(new_n783), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n399), .A2(new_n438), .ZN(new_n788));
  INV_X1    g602(.A(new_n579), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n599), .A2(new_n674), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n596), .A2(new_n788), .A3(new_n597), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n593), .B1(new_n348), .B2(new_n555), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n675), .A2(new_n655), .A3(new_n661), .ZN(new_n795));
  INV_X1    g609(.A(new_n584), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n683), .B1(new_n438), .B2(new_n603), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n561), .A2(new_n553), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n687), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n793), .A2(new_n684), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n775), .A2(new_n786), .A3(new_n787), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n781), .A2(new_n783), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n770), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT113), .B1(new_n769), .B2(new_n770), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n802), .B(new_n800), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n215), .A2(G952), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n758), .B2(new_n572), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n793), .A2(new_n799), .A3(KEYINPUT116), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n784), .A2(new_n812), .A3(new_n785), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT116), .B1(new_n793), .B2(new_n799), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n633), .A2(new_n637), .A3(new_n770), .ZN(new_n815));
  INV_X1    g629(.A(new_n684), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n787), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n811), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n753), .A2(new_n636), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n808), .A2(new_n810), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n750), .A2(new_n678), .A3(new_n755), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT48), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n823), .B(new_n825), .Z(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n824), .B2(KEYINPUT48), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n767), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(G952), .A2(G953), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n744), .B1(new_n828), .B2(new_n829), .ZN(G75));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n802), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n781), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n791), .B(KEYINPUT114), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n794), .A2(new_n687), .A3(new_n798), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n795), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n775), .A2(new_n787), .A3(new_n802), .A4(new_n800), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n224), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(G210), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n532), .A2(new_n533), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n516), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT55), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n215), .A2(G952), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G51));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n507), .B(KEYINPUT57), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT54), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(new_n820), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n857), .B2(new_n620), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT54), .B1(new_n840), .B2(new_n841), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n620), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(KEYINPUT120), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n840), .A2(new_n841), .A3(G902), .A4(new_n703), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT121), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n851), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n843), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n869), .A2(new_n395), .A3(new_n394), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n395), .B2(new_n394), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n870), .A2(new_n871), .A3(new_n851), .ZN(G60));
  NAND2_X1  g686(.A1(new_n568), .A2(new_n569), .ZN(new_n873));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT59), .Z(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n873), .B(new_n876), .C1(new_n859), .C2(new_n860), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n808), .B2(new_n820), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n867), .B(new_n877), .C1(new_n878), .C2(new_n873), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(G63));
  INV_X1    g694(.A(new_n842), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n228), .A2(new_n224), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n222), .A3(new_n221), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n591), .A3(new_n884), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n867), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(KEYINPUT61), .A3(new_n867), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(G66));
  AOI21_X1  g706(.A(new_n215), .B1(new_n441), .B2(G224), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n775), .A2(new_n794), .A3(new_n798), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n898), .B2(new_n215), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n846), .B1(G898), .B2(new_n215), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n899), .B(new_n900), .Z(G69));
  NAND2_X1  g715(.A1(G227), .A2(G900), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n724), .B1(new_n651), .B2(new_n677), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n711), .A2(new_n903), .A3(new_n726), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n782), .A2(new_n618), .A3(new_n687), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n736), .A3(new_n816), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n215), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n215), .A2(G900), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n387), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n302), .B(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(G953), .B(new_n902), .C1(new_n913), .C2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n902), .A2(G953), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n782), .A2(new_n615), .A3(new_n618), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n606), .A2(new_n674), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n348), .A2(new_n797), .A3(new_n925), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n727), .A2(new_n736), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n917), .B1(new_n927), .B2(G953), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n929), .ZN(G72));
  XNOR2_X1  g744(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n338), .A2(new_n224), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n898), .B2(new_n906), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n934), .A2(new_n303), .A3(new_n330), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n340), .B1(new_n326), .B2(new_n327), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n807), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n867), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n896), .A2(new_n927), .A3(new_n897), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n303), .B(new_n330), .C1(new_n939), .C2(new_n933), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n935), .A2(new_n938), .A3(new_n940), .ZN(G57));
endmodule


