

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U318 ( .A(n443), .B(n442), .ZN(n450) );
  XNOR2_X1 U319 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n442) );
  XNOR2_X1 U320 ( .A(n492), .B(n491), .ZN(n499) );
  XOR2_X1 U321 ( .A(n467), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U322 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n400) );
  XNOR2_X1 U323 ( .A(n416), .B(n400), .ZN(n401) );
  XNOR2_X1 U324 ( .A(n404), .B(n403), .ZN(n405) );
  INV_X1 U325 ( .A(KEYINPUT94), .ZN(n347) );
  NOR2_X1 U326 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U327 ( .A(n406), .B(n405), .ZN(n409) );
  XNOR2_X1 U328 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U329 ( .A(n350), .B(n349), .ZN(n353) );
  INV_X1 U330 ( .A(G162GAT), .ZN(n447) );
  XNOR2_X1 U331 ( .A(n355), .B(n354), .ZN(n516) );
  XNOR2_X1 U332 ( .A(n447), .B(KEYINPUT120), .ZN(n448) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(G1347GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n287) );
  XNOR2_X1 U335 ( .A(G99GAT), .B(G106GAT), .ZN(n286) );
  XNOR2_X1 U336 ( .A(n287), .B(n286), .ZN(n291) );
  XOR2_X1 U337 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n289) );
  XNOR2_X1 U338 ( .A(KEYINPUT11), .B(KEYINPUT66), .ZN(n288) );
  XNOR2_X1 U339 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U340 ( .A(n291), .B(n290), .Z(n301) );
  XOR2_X1 U341 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n293) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G29GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(KEYINPUT71), .B(n294), .Z(n394) );
  XOR2_X1 U345 ( .A(G162GAT), .B(KEYINPUT74), .Z(n296) );
  XNOR2_X1 U346 ( .A(G50GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n311) );
  XOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .Z(n337) );
  XOR2_X1 U349 ( .A(n311), .B(n337), .Z(n298) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n394), .B(n299), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(n302), .B(KEYINPUT9), .Z(n305) );
  XNOR2_X1 U355 ( .A(G92GAT), .B(G85GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n303), .B(KEYINPUT73), .ZN(n407) );
  XNOR2_X1 U357 ( .A(G190GAT), .B(n407), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n538) );
  XOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT87), .Z(n307) );
  XNOR2_X1 U360 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n370) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(G78GAT), .ZN(n308) );
  XOR2_X1 U363 ( .A(n308), .B(G148GAT), .Z(n398) );
  XNOR2_X1 U364 ( .A(n370), .B(n398), .ZN(n313) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT86), .Z(n310) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n351) );
  XNOR2_X1 U368 ( .A(n311), .B(n351), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U371 ( .A(KEYINPUT84), .B(KEYINPUT89), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U373 ( .A(n316), .B(KEYINPUT23), .Z(n318) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n382) );
  XNOR2_X1 U375 ( .A(n382), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U377 ( .A(KEYINPUT85), .B(KEYINPUT88), .Z(n320) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(G204GAT), .B(n321), .Z(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n467) );
  XOR2_X1 U383 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n327) );
  XNOR2_X1 U384 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U386 ( .A(n328), .B(G183GAT), .Z(n330) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(G176GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n355) );
  XOR2_X1 U389 ( .A(G127GAT), .B(KEYINPUT0), .Z(n332) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n359) );
  XOR2_X1 U392 ( .A(G99GAT), .B(G71GAT), .Z(n333) );
  XOR2_X1 U393 ( .A(G120GAT), .B(n333), .Z(n397) );
  XOR2_X1 U394 ( .A(n359), .B(n397), .Z(n341) );
  XOR2_X1 U395 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n335) );
  XNOR2_X1 U396 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U399 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U402 ( .A(n355), .B(n342), .Z(n526) );
  INV_X1 U403 ( .A(n526), .ZN(n518) );
  NOR2_X1 U404 ( .A1(n467), .A2(n518), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n343), .B(KEYINPUT26), .ZN(n562) );
  INV_X1 U406 ( .A(KEYINPUT114), .ZN(n445) );
  XNOR2_X1 U407 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n356) );
  XOR2_X1 U408 ( .A(G204GAT), .B(G64GAT), .Z(n402) );
  XOR2_X1 U409 ( .A(G92GAT), .B(G218GAT), .Z(n345) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G8GAT), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U412 ( .A(n402), .B(n346), .Z(n350) );
  NAND2_X1 U413 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n351), .B(KEYINPUT95), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n356), .B(n516), .ZN(n460) );
  XOR2_X1 U417 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U420 ( .A(n359), .B(KEYINPUT4), .Z(n361) );
  NAND2_X1 U421 ( .A1(G225GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n377) );
  XOR2_X1 U424 ( .A(G57GAT), .B(G148GAT), .Z(n365) );
  XNOR2_X1 U425 ( .A(G141GAT), .B(G120GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U427 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n367) );
  XNOR2_X1 U428 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U430 ( .A(n369), .B(n368), .Z(n375) );
  XOR2_X1 U431 ( .A(G85GAT), .B(n370), .Z(n372) );
  XNOR2_X1 U432 ( .A(G29GAT), .B(G162GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U434 ( .A(G134GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n514) );
  NAND2_X1 U437 ( .A1(n460), .A2(n514), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n378), .B(KEYINPUT97), .ZN(n468) );
  XOR2_X1 U439 ( .A(KEYINPUT67), .B(G197GAT), .Z(n380) );
  XNOR2_X1 U440 ( .A(G50GAT), .B(G43GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U442 ( .A(n381), .B(G113GAT), .Z(n384) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(n382), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U445 ( .A(G1GAT), .B(KEYINPUT72), .Z(n386) );
  XNOR2_X1 U446 ( .A(G15GAT), .B(G8GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n417) );
  XOR2_X1 U448 ( .A(n417), .B(KEYINPUT29), .Z(n388) );
  NAND2_X1 U449 ( .A1(G229GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n396) );
  XOR2_X1 U452 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U456 ( .A(n396), .B(n395), .Z(n501) );
  INV_X1 U457 ( .A(n501), .ZN(n564) );
  INV_X1 U458 ( .A(n397), .ZN(n399) );
  XOR2_X1 U459 ( .A(n399), .B(n398), .Z(n411) );
  XOR2_X1 U460 ( .A(KEYINPUT13), .B(G57GAT), .Z(n416) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n406) );
  NAND2_X1 U462 ( .A1(G230GAT), .A2(G233GAT), .ZN(n404) );
  INV_X1 U463 ( .A(KEYINPUT33), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n407), .B(KEYINPUT32), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n436) );
  XNOR2_X1 U467 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n436), .B(n412), .ZN(n552) );
  NOR2_X1 U469 ( .A1(n564), .A2(n552), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n413), .B(KEYINPUT46), .ZN(n431) );
  XOR2_X1 U471 ( .A(G78GAT), .B(G211GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(G22GAT), .B(G183GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n430) );
  XOR2_X1 U474 ( .A(n416), .B(G71GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(n417), .B(G127GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U477 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n421) );
  NAND2_X1 U478 ( .A1(G231GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n428) );
  XOR2_X1 U481 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n425) );
  XNOR2_X1 U482 ( .A(G155GAT), .B(G64GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n426), .B(KEYINPUT78), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n558) );
  INV_X1 U487 ( .A(n558), .ZN(n571) );
  NOR2_X1 U488 ( .A1(n431), .A2(n571), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n432), .B(KEYINPUT112), .ZN(n433) );
  AND2_X1 U490 ( .A1(n433), .A2(n538), .ZN(n435) );
  INV_X1 U491 ( .A(KEYINPUT47), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n441) );
  XNOR2_X1 U493 ( .A(KEYINPUT36), .B(n538), .ZN(n576) );
  NOR2_X1 U494 ( .A1(n576), .A2(n558), .ZN(n437) );
  XNOR2_X1 U495 ( .A(KEYINPUT45), .B(n437), .ZN(n438) );
  NAND2_X1 U496 ( .A1(n438), .A2(n564), .ZN(n439) );
  NOR2_X1 U497 ( .A1(n436), .A2(n439), .ZN(n440) );
  NOR2_X1 U498 ( .A1(n441), .A2(n440), .ZN(n443) );
  NAND2_X1 U499 ( .A1(n468), .A2(n450), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n528) );
  NAND2_X1 U501 ( .A1(n562), .A2(n528), .ZN(n446) );
  XNOR2_X1 U502 ( .A(KEYINPUT118), .B(n446), .ZN(n542) );
  NOR2_X1 U503 ( .A1(n538), .A2(n542), .ZN(n449) );
  XNOR2_X1 U504 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n452) );
  NAND2_X1 U505 ( .A1(n450), .A2(n516), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n561) );
  INV_X1 U507 ( .A(n514), .ZN(n560) );
  AND2_X1 U508 ( .A1(n467), .A2(n560), .ZN(n453) );
  NAND2_X1 U509 ( .A1(n561), .A2(n453), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n455), .A2(n518), .ZN(n557) );
  NOR2_X1 U512 ( .A1(n538), .A2(n557), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT58), .B(n456), .ZN(n458) );
  INV_X1 U514 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  NOR2_X1 U516 ( .A1(n564), .A2(n436), .ZN(n489) );
  NAND2_X1 U517 ( .A1(n538), .A2(n571), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n459), .Z(n475) );
  NAND2_X1 U519 ( .A1(n562), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT99), .B(n461), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n518), .A2(n516), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n467), .A2(n462), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n463), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n514), .A2(n466), .ZN(n473) );
  XOR2_X1 U526 ( .A(KEYINPUT82), .B(n518), .Z(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n527), .A2(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT98), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(n474), .Z(n486) );
  NAND2_X1 U531 ( .A1(n475), .A2(n486), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT101), .ZN(n502) );
  AND2_X1 U533 ( .A1(n489), .A2(n502), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n514), .A2(n483), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n516), .A2(n483), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U541 ( .A1(n483), .A2(n518), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n483), .A2(n527), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n576), .A2(n571), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(n488), .Z(n511) );
  NAND2_X1 U549 ( .A1(n489), .A2(n511), .ZN(n492) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n514), .A2(n499), .ZN(n494) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n516), .A2(n499), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n497) );
  NAND2_X1 U558 ( .A1(n499), .A2(n518), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U560 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n527), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n504) );
  NOR2_X1 U564 ( .A1(n501), .A2(n552), .ZN(n512) );
  AND2_X1 U565 ( .A1(n512), .A2(n502), .ZN(n508) );
  NAND2_X1 U566 ( .A1(n508), .A2(n514), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n516), .A2(n508), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n518), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n527), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(n513), .Z(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT109), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n521), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n525) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U587 ( .A1(n527), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n529) );
  NAND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n564), .A2(n537), .ZN(n530) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n552), .A2(n537), .ZN(n532) );
  XNOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NOR2_X1 U598 ( .A1(n558), .A2(n537), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n541), .Z(G1343GAT) );
  NOR2_X1 U606 ( .A1(n564), .A2(n542), .ZN(n543) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n552), .A2(n542), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n542), .A2(n558), .ZN(n548) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n564), .A2(n557), .ZN(n549) );
  XOR2_X1 U616 ( .A(G169GAT), .B(n549), .Z(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n552), .A2(n557), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  AND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n575) );
  NOR2_X1 U628 ( .A1(n575), .A2(n564), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n570) );
  INV_X1 U634 ( .A(n575), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n572), .A2(n436), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT126), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(n574), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

