//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT70), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G227gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G127gat), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G113gat), .ZN(new_n218));
  INV_X1    g017(.A(G113gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI211_X1 g029(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n230), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G169gat), .A3(G176gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n239), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n229), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(new_n232), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n240), .B1(new_n236), .B2(new_n255), .ZN(new_n256));
  NOR3_X1   g055(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n256), .A2(new_n257), .B1(new_n226), .B2(new_n227), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT27), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G183gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n260), .B1(new_n262), .B2(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n227), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n259), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND4_X1   g066(.A1(KEYINPUT28), .A2(new_n261), .A3(new_n263), .A4(new_n227), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n258), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n272), .B(new_n258), .C1(new_n267), .C2(new_n269), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n225), .B(new_n254), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT27), .B(G183gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n227), .B(new_n265), .C1(new_n276), .C2(new_n260), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n268), .B1(new_n277), .B2(new_n259), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n272), .B1(new_n278), .B2(new_n258), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n225), .B1(new_n281), .B2(new_n254), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n209), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n284));
  AOI21_X1  g083(.A(new_n206), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n209), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n254), .B1(new_n271), .B2(new_n273), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n216), .A2(new_n224), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n286), .B1(new_n289), .B2(new_n274), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(new_n293), .A3(KEYINPUT32), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n283), .B(KEYINPUT32), .C1(new_n284), .C2(new_n206), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n275), .A2(new_n282), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n286), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(new_n297), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT34), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n202), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT36), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n287), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  INV_X1    g117(.A(G218gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n315), .B1(new_n320), .B2(new_n316), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n278), .A2(new_n258), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n254), .A2(new_n324), .A3(new_n311), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n313), .A2(new_n314), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n242), .A2(new_n243), .B1(new_n252), .B2(new_n250), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n279), .B2(new_n280), .ZN(new_n328));
  INV_X1    g127(.A(new_n312), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n323), .B(new_n325), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n311), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n312), .B1(new_n327), .B2(new_n270), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(KEYINPUT37), .B(new_n326), .C1(new_n331), .C2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT73), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT83), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n326), .B1(new_n331), .B2(new_n334), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT37), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n335), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT38), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT2), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G155gat), .B(G162gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G141gat), .B(G148gat), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n351), .A2(KEYINPUT2), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n352), .B(new_n363), .C1(new_n366), .C2(new_n353), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(new_n367), .A3(KEYINPUT3), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n368), .A2(new_n288), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT75), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  AOI211_X1 g172(.A(new_n373), .B(KEYINPUT3), .C1(new_n358), .C2(new_n367), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n225), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT4), .B1(new_n225), .B2(new_n370), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n358), .A2(new_n367), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n288), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n225), .A2(new_n370), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n375), .A2(new_n378), .A3(KEYINPUT5), .A4(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  INV_X1    g194(.A(new_n393), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n396), .A3(new_n388), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n396), .A4(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n343), .A2(new_n339), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n339), .A2(KEYINPUT38), .ZN(new_n402));
  INV_X1    g201(.A(new_n323), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(new_n325), .C1(new_n328), .C2(new_n329), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT37), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n332), .B2(new_n333), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n344), .B2(new_n343), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n350), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n398), .A2(new_n400), .A3(new_n399), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n411), .A2(new_n408), .A3(KEYINPUT82), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n349), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n370), .A2(new_n371), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n373), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n372), .B2(new_n374), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n323), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n321), .B2(new_n322), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n371), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n425), .B2(new_n382), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n419), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(new_n417), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n403), .B1(new_n428), .B2(new_n420), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n403), .A2(KEYINPUT76), .A3(new_n420), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT76), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT3), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n370), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n423), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G22gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n427), .A2(new_n441), .A3(new_n434), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(KEYINPUT78), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n427), .A2(new_n434), .A3(new_n445), .A4(new_n441), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n446), .A3(new_n436), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n447), .A2(KEYINPUT79), .A3(new_n439), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT79), .B1(new_n447), .B2(new_n439), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n397), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  INV_X1    g251(.A(new_n378), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n368), .A2(new_n288), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n416), .B2(new_n417), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n452), .B(new_n381), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n393), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n459), .A3(new_n393), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n381), .B1(new_n453), .B2(new_n455), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n383), .A2(new_n384), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n462), .B(KEYINPUT39), .C1(new_n381), .C2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n451), .B1(new_n465), .B2(KEYINPUT40), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n400), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n339), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n343), .A2(new_n339), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n461), .A2(new_n464), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n472), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT81), .B1(new_n472), .B2(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n466), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n413), .A2(new_n450), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n306), .A2(new_n304), .A3(new_n298), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n202), .A3(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n398), .A2(new_n399), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  OAI221_X1 g282(.A(new_n443), .B1(new_n471), .B2(new_n483), .C1(new_n448), .C2(new_n449), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n310), .A2(new_n477), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n471), .A2(new_n483), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n450), .A2(new_n486), .A3(new_n479), .A4(new_n478), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n303), .A2(new_n307), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(new_n486), .A3(new_n450), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT85), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n485), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G232gat), .A2(G233gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT93), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT41), .ZN(new_n503));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT7), .ZN(new_n510));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  INV_X1    g310(.A(G85gat), .ZN(new_n512));
  INV_X1    g311(.A(G92gat), .ZN(new_n513));
  AOI22_X1  g312(.A1(KEYINPUT8), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G99gat), .B(G106gat), .Z(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n510), .A3(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(KEYINPUT96), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(G43gat), .A2(G50gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT88), .B(G50gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G43gat), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(G43gat), .A2(G50gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT15), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n531), .B1(new_n537), .B2(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(KEYINPUT87), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n538), .A2(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n536), .B1(new_n540), .B2(new_n534), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n524), .A2(new_n541), .B1(KEYINPUT41), .B2(new_n502), .ZN(new_n542));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT97), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n536), .B(KEYINPUT17), .C1(new_n534), .C2(new_n540), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n523), .A4(new_n522), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n542), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n545), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n508), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n508), .A2(new_n550), .A3(new_n551), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT98), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560));
  INV_X1    g359(.A(G71gat), .ZN(new_n561));
  INV_X1    g360(.A(G78gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n565), .A3(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n571), .A2(KEYINPUT10), .A3(new_n524), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n569), .A2(new_n570), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT92), .B1(new_n567), .B2(new_n568), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n520), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(new_n519), .A3(new_n517), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT10), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n558), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n571), .B2(new_n520), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n557), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n578), .A2(new_n581), .A3(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR3_X1    g389(.A1(new_n573), .A2(KEYINPUT21), .A3(new_n574), .ZN(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n212), .ZN(new_n594));
  XNOR2_X1  g393(.A(G15gat), .B(G22gat), .ZN(new_n595));
  INV_X1    g394(.A(G1gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT16), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(G1gat), .B2(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G8gat), .ZN(new_n600));
  INV_X1    g399(.A(G8gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n601), .C1(G1gat), .C2(new_n595), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n571), .B2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n594), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n593), .B(G127gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n605), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n605), .B2(new_n608), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n555), .B(new_n590), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n603), .B1(new_n541), .B2(new_n546), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n548), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n541), .A2(new_n603), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n617), .A2(KEYINPUT18), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(KEYINPUT13), .Z(new_n622));
  NOR2_X1   g421(.A1(new_n541), .A2(new_n603), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n541), .B(new_n603), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(KEYINPUT89), .A3(new_n622), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n618), .B1(new_n548), .B2(new_n616), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT18), .B1(new_n630), .B2(new_n620), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT11), .B(G169gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n620), .A3(new_n619), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT18), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT90), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n638), .B1(new_n631), .B2(KEYINPUT90), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(KEYINPUT91), .A3(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n640), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n615), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n499), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n483), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n471), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n601), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n658), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n655), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n655), .A2(new_n657), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(KEYINPUT100), .B(new_n661), .C1(new_n655), .C2(new_n657), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(new_n652), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n308), .A2(new_n309), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT36), .B1(new_n480), .B2(new_n202), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G15gat), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n480), .A2(G15gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n666), .B2(new_n671), .ZN(G1326gat));
  INV_X1    g471(.A(new_n450), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(G29gat), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n555), .A2(KEYINPUT103), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n555), .A2(KEYINPUT103), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n485), .A2(KEYINPUT101), .B1(new_n489), .B2(new_n493), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n685), .A3(new_n477), .A4(new_n484), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n553), .A2(new_n554), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n496), .A2(new_n498), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(KEYINPUT44), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n613), .A2(new_n614), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n650), .A3(new_n589), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n677), .B1(new_n695), .B2(new_n483), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n496), .A2(new_n498), .A3(new_n688), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n483), .A2(new_n677), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n696), .B2(new_n700), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1328gat));
  INV_X1    g503(.A(new_n695), .ZN(new_n705));
  INV_X1    g504(.A(new_n471), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n697), .A2(G36gat), .A3(new_n706), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n669), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G43gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n480), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n697), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n713), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g521(.A(new_n712), .B(new_n720), .C1(new_n715), .C2(G43gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n690), .A2(new_n450), .A3(new_n694), .ZN(new_n726));
  INV_X1    g525(.A(new_n527), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n673), .A2(new_n727), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n697), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n730), .B2(new_n697), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n726), .B2(new_n727), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(new_n733), .A3(KEYINPUT48), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  OAI221_X1 g534(.A(new_n732), .B1(new_n725), .B2(new_n735), .C1(new_n726), .C2(new_n727), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n734), .A2(new_n736), .ZN(G1331gat));
  NAND4_X1  g536(.A1(new_n692), .A2(new_n650), .A3(new_n555), .A4(new_n589), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n684), .B2(new_n686), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n483), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n471), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  AOI21_X1  g544(.A(new_n561), .B1(new_n739), .B2(new_n714), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n480), .A2(G71gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n739), .A2(new_n673), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  INV_X1    g550(.A(new_n690), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n644), .A2(KEYINPUT91), .A3(new_n645), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT91), .B1(new_n644), .B2(new_n645), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n753), .A2(new_n754), .B1(new_n639), .B2(new_n632), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n692), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n589), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n482), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n684), .A2(new_n686), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n692), .A2(new_n755), .A3(new_n555), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n512), .A3(new_n483), .A4(new_n589), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(new_n764), .ZN(G1336gat));
  NAND4_X1  g564(.A1(new_n752), .A2(new_n471), .A3(new_n589), .A4(new_n756), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n706), .A2(G92gat), .A3(new_n590), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT108), .B1(new_n759), .B2(new_n760), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT51), .Z(new_n772));
  AOI22_X1  g571(.A1(new_n772), .A2(new_n768), .B1(new_n766), .B2(G92gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n757), .B2(new_n669), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n480), .A2(G99gat), .A3(new_n590), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1338gat));
  OR3_X1    g578(.A1(new_n450), .A2(G106gat), .A3(new_n590), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n752), .A2(new_n673), .A3(new_n589), .A4(new_n756), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT109), .B(G106gat), .Z(new_n783));
  AOI22_X1  g582(.A1(new_n772), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n761), .B2(new_n762), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n782), .A2(new_n783), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n784), .A2(new_n785), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  NOR2_X1   g591(.A1(new_n615), .A2(new_n755), .ZN(new_n793));
  INV_X1    g592(.A(new_n636), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n627), .A2(new_n622), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT113), .Z(new_n796));
  OR2_X1    g595(.A1(new_n630), .A2(new_n620), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n648), .B2(new_n649), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n571), .A2(new_n524), .A3(KEYINPUT10), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n557), .B(new_n800), .C1(new_n580), .C2(KEYINPUT10), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n578), .A2(new_n801), .A3(KEYINPUT54), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n578), .A2(new_n801), .A3(KEYINPUT112), .A4(KEYINPUT54), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n806), .B(new_n558), .C1(new_n572), .C2(new_n577), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n586), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n588), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n586), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n803), .B2(new_n802), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n812), .B2(new_n805), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n681), .A2(new_n799), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n797), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n636), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n589), .C1(new_n754), .C2(new_n753), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n588), .A3(new_n809), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT114), .B(new_n818), .C1(new_n822), .C2(new_n650), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n680), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n809), .A2(new_n588), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n755), .A3(new_n821), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT114), .B1(new_n826), .B2(new_n818), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n815), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n793), .B1(new_n828), .B2(new_n691), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n673), .A2(new_n480), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n829), .A2(new_n482), .A3(new_n471), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n755), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT115), .B1(new_n829), .B2(new_n673), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n490), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n471), .A2(new_n482), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n828), .A2(new_n691), .ZN(new_n837));
  INV_X1    g636(.A(new_n793), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n450), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n650), .A2(new_n219), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n833), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  AOI21_X1  g644(.A(G120gat), .B1(new_n832), .B2(new_n589), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n590), .A2(new_n217), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n843), .B2(new_n847), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n842), .B2(new_n691), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n212), .A3(new_n692), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n210), .A3(new_n688), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT56), .Z(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n842), .B2(new_n555), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n669), .A2(new_n836), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n818), .B1(new_n822), .B2(new_n650), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n555), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n815), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n793), .B1(new_n860), .B2(new_n691), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n673), .A2(KEYINPUT57), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n450), .B1(new_n837), .B2(new_n838), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n857), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n650), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n829), .A2(new_n482), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n669), .A2(new_n673), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n471), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(G141gat), .A3(new_n650), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT58), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(new_n857), .C1(new_n866), .C2(new_n868), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n755), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n875), .B1(KEYINPUT118), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n877), .B1(new_n882), .B2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(new_n874), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n361), .A3(new_n589), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G148gat), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n878), .A2(new_n880), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n589), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n814), .A2(new_n688), .A3(new_n799), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n814), .A2(new_n755), .B1(new_n589), .B2(new_n799), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n688), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n793), .B1(new_n895), .B2(new_n691), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(new_n450), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n867), .A2(KEYINPUT57), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR4_X1   g698(.A1(new_n829), .A2(KEYINPUT119), .A3(new_n892), .A4(new_n450), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n589), .B(new_n857), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n888), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n887), .B1(new_n891), .B2(new_n902), .ZN(G1345gat));
  AOI21_X1  g702(.A(KEYINPUT120), .B1(new_n886), .B2(new_n692), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n874), .A2(new_n905), .A3(new_n691), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n904), .A2(G155gat), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n692), .A2(G155gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n890), .B2(new_n908), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n878), .A2(new_n681), .A3(new_n880), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n878), .A2(new_n912), .A3(new_n681), .A4(new_n880), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(G162gat), .A3(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n874), .A2(G162gat), .A3(new_n555), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT121), .Z(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n706), .A2(new_n483), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n841), .A2(new_n834), .A3(new_n490), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n650), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n839), .A2(new_n482), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(new_n706), .A3(new_n831), .ZN(new_n922));
  INV_X1    g721(.A(G169gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n755), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT123), .Z(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n919), .B2(new_n590), .ZN(new_n927));
  INV_X1    g726(.A(G176gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n922), .A2(new_n928), .A3(new_n589), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1349gat));
  NAND3_X1  g729(.A1(new_n922), .A2(new_n276), .A3(new_n692), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n919), .B2(new_n691), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G183gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n691), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT60), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n938), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n227), .A3(new_n681), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n919), .A2(new_n555), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(G190gat), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n942), .B2(G190gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n921), .A2(new_n706), .A3(new_n872), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n755), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n669), .A2(new_n918), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT114), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n858), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n680), .A3(new_n823), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n692), .B1(new_n953), .B2(new_n815), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT57), .B(new_n673), .C1(new_n954), .C2(new_n793), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n688), .B1(new_n826), .B2(new_n818), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n814), .A2(new_n688), .A3(new_n799), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n691), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n450), .B1(new_n958), .B2(new_n838), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n898), .B1(new_n959), .B2(KEYINPUT57), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n839), .A2(new_n898), .A3(KEYINPUT57), .A4(new_n673), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n950), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n755), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n949), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n966), .A3(new_n589), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  AND2_X1   g767(.A1(new_n963), .A2(new_n589), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n966), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n948), .A2(new_n318), .A3(new_n692), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n972));
  AOI211_X1 g771(.A(new_n972), .B(new_n318), .C1(new_n963), .C2(new_n692), .ZN(new_n973));
  INV_X1    g772(.A(new_n950), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n692), .B(new_n974), .C1(new_n899), .C2(new_n900), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n971), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n979), .B(new_n971), .C1(new_n973), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1354gat));
  AOI21_X1  g780(.A(new_n319), .B1(new_n963), .B2(new_n688), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n680), .A2(G218gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n948), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n984), .B(new_n985), .ZN(G1355gat));
endmodule


