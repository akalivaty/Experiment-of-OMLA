

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U555 ( .A1(n735), .A2(n734), .ZN(n733) );
  NOR2_X1 U556 ( .A1(n764), .A2(n933), .ZN(n724) );
  AND2_X1 U557 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X4 U558 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  NOR2_X1 U559 ( .A1(G1384), .A2(n709), .ZN(n722) );
  NOR2_X1 U560 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U561 ( .A1(n885), .A2(G137), .ZN(n528) );
  XOR2_X1 U562 ( .A(KEYINPUT14), .B(n571), .Z(n523) );
  INV_X1 U563 ( .A(n809), .ZN(n790) );
  NAND2_X1 U564 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U565 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U566 ( .A(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U567 ( .A1(G651), .A2(n646), .ZN(n651) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n538), .Z(n649) );
  NOR2_X1 U569 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U570 ( .A(KEYINPUT65), .ZN(n536) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U572 ( .A(n525), .B(n524), .ZN(n885) );
  XOR2_X2 U573 ( .A(KEYINPUT66), .B(n526), .Z(n882) );
  NAND2_X1 U574 ( .A1(n882), .A2(G113), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n529), .B(KEYINPUT67), .ZN(n535) );
  INV_X1 U577 ( .A(G2105), .ZN(n530) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n530), .ZN(n881) );
  AND2_X1 U579 ( .A1(G125), .A2(n881), .ZN(n533) );
  AND2_X1 U580 ( .A1(n530), .A2(G2104), .ZN(n886) );
  NAND2_X1 U581 ( .A1(G101), .A2(n886), .ZN(n531) );
  XNOR2_X1 U582 ( .A(KEYINPUT23), .B(n531), .ZN(n532) );
  NOR2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X2 U584 ( .A(n537), .B(n536), .ZN(G160) );
  XOR2_X1 U585 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  NAND2_X1 U586 ( .A1(G53), .A2(n651), .ZN(n540) );
  INV_X1 U587 ( .A(G651), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G543), .A2(n541), .ZN(n538) );
  NAND2_X1 U589 ( .A1(G65), .A2(n649), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U591 ( .A1(G91), .A2(n652), .ZN(n543) );
  NOR2_X1 U592 ( .A1(n646), .A2(n541), .ZN(n655) );
  NAND2_X1 U593 ( .A1(G78), .A2(n655), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U595 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U596 ( .A(n546), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U597 ( .A1(G52), .A2(n651), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G64), .A2(n649), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U600 ( .A(KEYINPUT69), .B(n549), .Z(n555) );
  NAND2_X1 U601 ( .A1(n655), .A2(G77), .ZN(n550) );
  XNOR2_X1 U602 ( .A(n550), .B(KEYINPUT70), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G90), .A2(n652), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U606 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U607 ( .A1(G138), .A2(n885), .ZN(n557) );
  NAND2_X1 U608 ( .A1(G102), .A2(n886), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT91), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G114), .A2(n882), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U613 ( .A1(G126), .A2(n881), .ZN(n561) );
  XOR2_X1 U614 ( .A(KEYINPUT90), .B(n561), .Z(n562) );
  XNOR2_X1 U615 ( .A(n564), .B(KEYINPUT92), .ZN(n709) );
  BUF_X1 U616 ( .A(n709), .Z(G164) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G860), .ZN(n610) );
  NAND2_X1 U619 ( .A1(n652), .A2(G81), .ZN(n565) );
  XNOR2_X1 U620 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G68), .A2(n655), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U623 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U624 ( .A1(G43), .A2(n651), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n649), .A2(G56), .ZN(n571) );
  NOR2_X1 U627 ( .A1(n572), .A2(n523), .ZN(n573) );
  XOR2_X2 U628 ( .A(KEYINPUT74), .B(n573), .Z(n949) );
  OR2_X1 U629 ( .A1(n610), .A2(n949), .ZN(G153) );
  INV_X1 U630 ( .A(G120), .ZN(G236) );
  INV_X1 U631 ( .A(G69), .ZN(G235) );
  INV_X1 U632 ( .A(G108), .ZN(G238) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G88), .A2(n652), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G75), .A2(n655), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G50), .A2(n651), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G62), .A2(n649), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(G166) );
  NAND2_X1 U642 ( .A1(G51), .A2(n651), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G63), .A2(n649), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT6), .B(n582), .ZN(n590) );
  NAND2_X1 U646 ( .A1(G89), .A2(n652), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT4), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT76), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G76), .A2(n655), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT5), .B(n587), .ZN(n588) );
  XNOR2_X1 U652 ( .A(KEYINPUT77), .B(n588), .ZN(n589) );
  NOR2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT7), .B(n591), .Z(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(KEYINPUT72), .ZN(n593) );
  XNOR2_X1 U658 ( .A(KEYINPUT10), .B(n593), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n837) );
  NAND2_X1 U660 ( .A1(n837), .A2(G567), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT73), .ZN(n595) );
  XNOR2_X1 U662 ( .A(KEYINPUT11), .B(n595), .ZN(G234) );
  NAND2_X1 U663 ( .A1(G868), .A2(G171), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G54), .A2(n651), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G66), .A2(n649), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G92), .A2(n652), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G79), .A2(n655), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT15), .ZN(n734) );
  INV_X1 U672 ( .A(n734), .ZN(n955) );
  INV_X1 U673 ( .A(G868), .ZN(n670) );
  NAND2_X1 U674 ( .A1(n955), .A2(n670), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT75), .ZN(G284) );
  NOR2_X1 U677 ( .A1(G286), .A2(n670), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT78), .B(n606), .Z(n608) );
  INV_X1 U679 ( .A(G299), .ZN(n958) );
  NAND2_X1 U680 ( .A1(n958), .A2(n670), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT79), .B(n609), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n611), .A2(n955), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(n949), .A2(G868), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G868), .A2(n955), .ZN(n613) );
  NOR2_X1 U688 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(G282) );
  XOR2_X1 U690 ( .A(G2100), .B(KEYINPUT80), .Z(n624) );
  NAND2_X1 U691 ( .A1(G123), .A2(n881), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n886), .A2(G99), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G135), .A2(n885), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G111), .A2(n882), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n1010) );
  XNOR2_X1 U699 ( .A(n1010), .B(G2096), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G55), .A2(n651), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G67), .A2(n649), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G93), .A2(n652), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G80), .A2(n655), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n669) );
  NAND2_X1 U708 ( .A1(G559), .A2(n955), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n631), .B(KEYINPUT81), .ZN(n667) );
  XOR2_X1 U710 ( .A(n667), .B(n949), .Z(n632) );
  NOR2_X1 U711 ( .A1(G860), .A2(n632), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT82), .B(n633), .Z(n634) );
  XOR2_X1 U713 ( .A(n669), .B(n634), .Z(G145) );
  NAND2_X1 U714 ( .A1(G85), .A2(n652), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G72), .A2(n655), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G47), .A2(n651), .ZN(n637) );
  XOR2_X1 U718 ( .A(KEYINPUT68), .B(n637), .Z(n638) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n649), .A2(G60), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G49), .A2(n651), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n649), .A2(n644), .ZN(n645) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n645), .Z(n648) );
  NAND2_X1 U727 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G61), .A2(n649), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n650), .B(KEYINPUT84), .ZN(n660) );
  NAND2_X1 U731 ( .A1(G48), .A2(n651), .ZN(n654) );
  NAND2_X1 U732 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(G305) );
  XNOR2_X1 U738 ( .A(n669), .B(G290), .ZN(n666) );
  XNOR2_X1 U739 ( .A(G288), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n949), .B(G166), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n958), .B(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n903) );
  XNOR2_X1 U745 ( .A(n667), .B(n903), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U749 ( .A(KEYINPUT85), .B(n673), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U754 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U758 ( .A1(G218), .A2(n679), .ZN(n680) );
  XNOR2_X1 U759 ( .A(KEYINPUT86), .B(n680), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(G96), .ZN(n842) );
  AND2_X1 U761 ( .A1(G2106), .A2(n842), .ZN(n687) );
  NOR2_X1 U762 ( .A1(G235), .A2(G236), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n682), .B(KEYINPUT87), .ZN(n683) );
  NOR2_X1 U764 ( .A1(G238), .A2(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G57), .A2(n684), .ZN(n841) );
  NAND2_X1 U766 ( .A1(G567), .A2(n841), .ZN(n685) );
  XOR2_X1 U767 ( .A(KEYINPUT88), .B(n685), .Z(n686) );
  NOR2_X1 U768 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U772 ( .A(KEYINPUT89), .B(n690), .Z(n840) );
  NAND2_X1 U773 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  NAND2_X1 U775 ( .A1(G141), .A2(n885), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G129), .A2(n881), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n886), .A2(G105), .ZN(n693) );
  XOR2_X1 U779 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U781 ( .A1(G117), .A2(n882), .ZN(n696) );
  NAND2_X1 U782 ( .A1(n697), .A2(n696), .ZN(n878) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n878), .ZN(n698) );
  XNOR2_X1 U784 ( .A(n698), .B(KEYINPUT95), .ZN(n708) );
  NAND2_X1 U785 ( .A1(G131), .A2(n885), .ZN(n700) );
  NAND2_X1 U786 ( .A1(G95), .A2(n886), .ZN(n699) );
  NAND2_X1 U787 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U788 ( .A(KEYINPUT94), .B(n701), .Z(n703) );
  NAND2_X1 U789 ( .A1(G107), .A2(n882), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G119), .A2(n881), .ZN(n704) );
  XNOR2_X1 U792 ( .A(KEYINPUT93), .B(n704), .ZN(n705) );
  OR2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n870) );
  AND2_X1 U794 ( .A1(G1991), .A2(n870), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n1007) );
  NOR2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n832) );
  INV_X1 U797 ( .A(n832), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n1007), .A2(n710), .ZN(n822) );
  INV_X1 U799 ( .A(n822), .ZN(n720) );
  NAND2_X1 U800 ( .A1(G140), .A2(n885), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G104), .A2(n886), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U803 ( .A(KEYINPUT34), .B(n713), .ZN(n718) );
  NAND2_X1 U804 ( .A1(G128), .A2(n881), .ZN(n715) );
  NAND2_X1 U805 ( .A1(G116), .A2(n882), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U807 ( .A(KEYINPUT35), .B(n716), .Z(n717) );
  NOR2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT36), .B(n719), .ZN(n899) );
  XNOR2_X1 U810 ( .A(G2067), .B(KEYINPUT37), .ZN(n829) );
  NOR2_X1 U811 ( .A1(n899), .A2(n829), .ZN(n1009) );
  NAND2_X1 U812 ( .A1(n832), .A2(n1009), .ZN(n827) );
  NAND2_X1 U813 ( .A1(n720), .A2(n827), .ZN(n817) );
  INV_X1 U814 ( .A(n721), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n764) );
  INV_X1 U816 ( .A(G1996), .ZN(n933) );
  XOR2_X1 U817 ( .A(KEYINPUT26), .B(n724), .Z(n726) );
  NAND2_X1 U818 ( .A1(n764), .A2(G1341), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X2 U820 ( .A1(n727), .A2(n949), .ZN(n728) );
  XOR2_X1 U821 ( .A(n728), .B(KEYINPUT64), .Z(n735) );
  AND2_X1 U822 ( .A1(n764), .A2(G1348), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT99), .ZN(n731) );
  INV_X1 U824 ( .A(n764), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n750), .A2(G2067), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n750), .A2(G2072), .ZN(n738) );
  XNOR2_X1 U831 ( .A(n738), .B(KEYINPUT27), .ZN(n740) );
  INV_X1 U832 ( .A(G1956), .ZN(n974) );
  NOR2_X1 U833 ( .A1(n974), .A2(n750), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n743), .A2(n958), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n743), .A2(n958), .ZN(n745) );
  XOR2_X1 U838 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n744) );
  XNOR2_X1 U839 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U841 ( .A(n748), .B(KEYINPUT29), .Z(n755) );
  NOR2_X1 U842 ( .A1(n750), .A2(G1961), .ZN(n749) );
  XOR2_X1 U843 ( .A(KEYINPUT96), .B(n749), .Z(n752) );
  XNOR2_X1 U844 ( .A(G2078), .B(KEYINPUT25), .ZN(n932) );
  NAND2_X1 U845 ( .A1(n750), .A2(n932), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n756) );
  AND2_X1 U847 ( .A1(n756), .A2(G171), .ZN(n753) );
  XNOR2_X1 U848 ( .A(KEYINPUT97), .B(n753), .ZN(n754) );
  NAND2_X1 U849 ( .A1(n755), .A2(n754), .ZN(n775) );
  NOR2_X1 U850 ( .A1(G171), .A2(n756), .ZN(n757) );
  XNOR2_X1 U851 ( .A(n757), .B(KEYINPUT100), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G8), .A2(n764), .ZN(n809) );
  NOR2_X1 U853 ( .A1(G1966), .A2(n809), .ZN(n781) );
  NOR2_X1 U854 ( .A1(G2084), .A2(n764), .ZN(n777) );
  NOR2_X1 U855 ( .A1(n781), .A2(n777), .ZN(n758) );
  NAND2_X1 U856 ( .A1(G8), .A2(n758), .ZN(n759) );
  XNOR2_X1 U857 ( .A(KEYINPUT30), .B(n759), .ZN(n760) );
  NOR2_X1 U858 ( .A1(n760), .A2(G168), .ZN(n761) );
  NOR2_X1 U859 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U860 ( .A(KEYINPUT31), .B(n763), .Z(n776) );
  NOR2_X1 U861 ( .A1(G1971), .A2(n809), .ZN(n766) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n764), .ZN(n765) );
  NOR2_X1 U863 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U864 ( .A1(n767), .A2(G303), .ZN(n769) );
  AND2_X1 U865 ( .A1(n776), .A2(n769), .ZN(n768) );
  NAND2_X1 U866 ( .A1(n775), .A2(n768), .ZN(n773) );
  INV_X1 U867 ( .A(n769), .ZN(n770) );
  OR2_X1 U868 ( .A1(n770), .A2(G286), .ZN(n771) );
  AND2_X1 U869 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U871 ( .A(KEYINPUT32), .B(n774), .Z(n783) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U873 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X2 U876 ( .A1(n783), .A2(n782), .ZN(n794) );
  INV_X1 U877 ( .A(G1971), .ZN(n988) );
  NAND2_X1 U878 ( .A1(G166), .A2(n988), .ZN(n784) );
  OR2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n784), .A2(n785), .ZN(n964) );
  NOR2_X1 U881 ( .A1(n794), .A2(n964), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n965) );
  INV_X1 U883 ( .A(KEYINPUT33), .ZN(n798) );
  OR2_X1 U884 ( .A1(n809), .A2(n785), .ZN(n786) );
  NOR2_X1 U885 ( .A1(n798), .A2(n786), .ZN(n787) );
  XNOR2_X1 U886 ( .A(n787), .B(KEYINPUT101), .ZN(n797) );
  AND2_X1 U887 ( .A1(n965), .A2(n797), .ZN(n789) );
  XNOR2_X1 U888 ( .A(G1981), .B(G305), .ZN(n951) );
  INV_X1 U889 ( .A(n951), .ZN(n788) );
  AND2_X1 U890 ( .A1(n789), .A2(n788), .ZN(n791) );
  OR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n814) );
  INV_X1 U892 ( .A(n794), .ZN(n807) );
  NOR2_X1 U893 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U894 ( .A1(G8), .A2(n795), .ZN(n796) );
  XNOR2_X1 U895 ( .A(n796), .B(KEYINPUT102), .ZN(n805) );
  INV_X1 U896 ( .A(n797), .ZN(n799) );
  OR2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n951), .A2(n800), .ZN(n804) );
  NOR2_X1 U899 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U900 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  NOR2_X1 U901 ( .A1(n809), .A2(n802), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U903 ( .A1(n805), .A2(n808), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n812) );
  INV_X1 U905 ( .A(n808), .ZN(n810) );
  OR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT103), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n819) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n960) );
  NAND2_X1 U912 ( .A1(n960), .A2(n832), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n835) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n878), .ZN(n1020) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n870), .ZN(n1011) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n1011), .A2(n820), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT104), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n1020), .A2(n824), .ZN(n826) );
  XOR2_X1 U921 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n825) );
  XNOR2_X1 U922 ( .A(n826), .B(n825), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n899), .A2(n829), .ZN(n1025) );
  NAND2_X1 U925 ( .A1(n830), .A2(n1025), .ZN(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT106), .B(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n836), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(G2100), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2090), .B(KEYINPUT110), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(G2678), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2096), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1976), .B(G1956), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(G1971), .B(G1986), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U956 ( .A(KEYINPUT111), .B(G2474), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U958 ( .A(G1981), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G100), .A2(n886), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G112), .A2(n882), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(n864), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G124), .A2(n881), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n885), .A2(G136), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(n870), .B(G162), .Z(n898) );
  XNOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G139), .A2(n885), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G103), .A2(n886), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G127), .A2(n881), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G115), .A2(n882), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n1015) );
  XNOR2_X1 U979 ( .A(n878), .B(n1015), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n894) );
  NAND2_X1 U981 ( .A1(G130), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n892) );
  NAND2_X1 U984 ( .A1(G142), .A2(n885), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G106), .A2(n886), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(n889), .ZN(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT45), .B(n890), .ZN(n891) );
  NOR2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U991 ( .A(G164), .B(n1010), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n901) );
  XOR2_X1 U994 ( .A(n899), .B(G160), .Z(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT114), .B(n903), .Z(n905) );
  XNOR2_X1 U998 ( .A(n955), .B(G286), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(G171), .B(n906), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n907), .ZN(G397) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2446), .ZN(n917) );
  XOR2_X1 U1003 ( .A(G2430), .B(KEYINPUT108), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G2451), .B(G2443), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1006 ( .A(G2427), .B(KEYINPUT107), .Z(n911) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2435), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n918), .A2(G14), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G57), .ZN(G237) );
  INV_X1 U1022 ( .A(n924), .ZN(G401) );
  XOR2_X1 U1023 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1036) );
  XOR2_X1 U1024 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1030) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(G2090), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(G35), .ZN(n944) );
  XNOR2_X1 U1027 ( .A(G2084), .B(KEYINPUT54), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(n926), .B(G34), .ZN(n942) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(G2072), .B(G33), .ZN(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(n929), .B(KEYINPUT120), .ZN(n931) );
  XOR2_X1 U1033 ( .A(G1991), .B(G25), .Z(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n932), .B(G27), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n933), .B(G32), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(n936), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n937), .A2(G28), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(n940), .B(KEYINPUT53), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n1030), .B(n945), .ZN(n947) );
  INV_X1 U1045 ( .A(G29), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n948), .ZN(n1004) );
  XNOR2_X1 U1048 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XNOR2_X1 U1049 ( .A(n949), .B(G1341), .ZN(n954) );
  XOR2_X1 U1050 ( .A(G1966), .B(G168), .Z(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT57), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n971) );
  XNOR2_X1 U1054 ( .A(G1348), .B(n955), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G171), .B(G1961), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(n958), .B(G1956), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(G166), .A2(n988), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT122), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1002) );
  INV_X1 U1067 ( .A(G16), .ZN(n1000) );
  XOR2_X1 U1068 ( .A(G1961), .B(G5), .Z(n987) );
  XNOR2_X1 U1069 ( .A(G20), .B(n974), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n975), .B(KEYINPUT123), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G6), .B(G1981), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(n980), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n981), .B(G4), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(n984), .B(KEYINPUT125), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT60), .B(n985), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n997) );
  XOR2_X1 U1082 ( .A(G1966), .B(G21), .Z(n995) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n990) );
  XNOR2_X1 U1084 ( .A(n988), .B(G22), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(KEYINPUT58), .B(n993), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT61), .B(n998), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1034) );
  XOR2_X1 U1095 ( .A(G160), .B(G2084), .Z(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT115), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT116), .B(n1014), .ZN(n1028) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1015), .Z(n1017) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1018), .Z(n1024) );
  XOR2_X1 U1106 ( .A(G2090), .B(G162), .Z(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(KEYINPUT117), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT51), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(KEYINPUT52), .B(n1029), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(G29), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(n1036), .B(n1035), .ZN(G311) );
  XNOR2_X1 U1118 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1119 ( .A(G171), .ZN(G301) );
endmodule

