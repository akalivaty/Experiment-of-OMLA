//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n453), .A2(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT71), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n474), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n477), .B2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n474), .A2(new_n477), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G124), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n489), .A2(new_n465), .A3(new_n467), .A4(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n477), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n477), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G62), .A3(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(new_n511), .B1(new_n508), .B2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n505), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n500), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT7), .Z(new_n521));
  AND3_X1   g096(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n513), .ZN(new_n523));
  AOI211_X1 g098(.A(new_n521), .B(new_n522), .C1(G89), .C2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n512), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n500), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n510), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G52), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(G90), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n504), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n526), .A2(G43), .B1(G651), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n523), .A2(G81), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(new_n523), .A2(G91), .ZN(new_n547));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n504), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n512), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n547), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(G299));
  INV_X1    g131(.A(G168), .ZN(G286));
  INV_X1    g132(.A(G166), .ZN(G303));
  NAND2_X1  g133(.A1(new_n526), .A2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n523), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  AOI22_X1  g137(.A1(new_n526), .A2(G48), .B1(new_n523), .B2(G86), .ZN(new_n563));
  INV_X1    g138(.A(G61), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n504), .A2(KEYINPUT74), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT74), .B1(new_n504), .B2(new_n564), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n563), .A2(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n510), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT75), .Z(new_n573));
  AOI22_X1  g148(.A1(new_n526), .A2(G47), .B1(new_n523), .B2(G85), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n523), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT76), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT77), .B(G66), .Z(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n504), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT78), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(G54), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G284));
  XNOR2_X1  g163(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  XNOR2_X1  g165(.A(G299), .B(KEYINPUT80), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(G868), .B2(new_n591), .ZN(G297));
  OAI21_X1  g167(.A(new_n590), .B1(G868), .B2(new_n591), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n587), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g174(.A1(new_n481), .A2(G135), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n486), .A2(G123), .ZN(new_n603));
  OR2_X1    g178(.A1(G99), .A2(G2105), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n604), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n481), .A2(KEYINPUT82), .A3(G135), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n602), .A2(new_n603), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2096), .Z(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n466), .A2(new_n464), .A3(G2105), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT13), .B(G2100), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(G156));
  XOR2_X1   g189(.A(KEYINPUT15), .B(G2435), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2438), .ZN(new_n616));
  XOR2_X1   g191(.A(G2427), .B(G2430), .Z(new_n617));
  OAI21_X1  g192(.A(KEYINPUT14), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT83), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n616), .A2(new_n617), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT85), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2443), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G14), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(G401));
  XNOR2_X1  g207(.A(G2084), .B(G2090), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT86), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2072), .B(G2078), .ZN(new_n635));
  XOR2_X1   g210(.A(G2067), .B(G2678), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT87), .Z(new_n639));
  XOR2_X1   g214(.A(new_n635), .B(KEYINPUT17), .Z(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n636), .ZN(new_n641));
  INV_X1    g216(.A(new_n634), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n642), .A2(new_n640), .A3(new_n636), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n635), .A3(new_n637), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT18), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n641), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G227));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT88), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT19), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n653), .A2(new_n656), .A3(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G1981), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  AOI22_X1  g243(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n669), .A2(new_n477), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT93), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n481), .A2(G139), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT25), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(G33), .B(new_n675), .S(G29), .Z(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2072), .Z(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G27), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G164), .B2(new_n678), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2078), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(G168), .A2(G16), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G21), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(KEYINPUT98), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(KEYINPUT98), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT99), .B(G1966), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT100), .B(KEYINPUT31), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G11), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(G28), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(G28), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n693), .A3(new_n678), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n690), .B(new_n694), .C1(new_n607), .C2(new_n678), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT101), .Z(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n686), .B2(new_n687), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(new_n678), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n479), .B2(new_n678), .ZN(new_n701));
  INV_X1    g276(.A(G2084), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n678), .A2(G32), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n477), .A2(G105), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT95), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n481), .A2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n486), .A2(G129), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n704), .B1(new_n714), .B2(new_n678), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT97), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n688), .A2(new_n697), .A3(new_n703), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G171), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G5), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(KEYINPUT102), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n701), .A2(new_n702), .ZN(new_n726));
  NOR4_X1   g301(.A1(new_n682), .A2(new_n719), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT103), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n731), .A2(KEYINPUT23), .A3(G20), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n733));
  INV_X1    g308(.A(G20), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G299), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n735), .C1(new_n736), .C2(new_n731), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1956), .Z(new_n738));
  AND2_X1   g313(.A1(new_n678), .A2(G26), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n481), .A2(G140), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT92), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n486), .A2(G128), .ZN(new_n742));
  NOR2_X1   g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(new_n477), .B2(G116), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  MUX2_X1   g321(.A(new_n739), .B(new_n746), .S(KEYINPUT28), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2067), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n729), .A2(new_n730), .A3(new_n738), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT29), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n756));
  MUX2_X1   g331(.A(G6), .B(G305), .S(G16), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1981), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n731), .A2(G23), .ZN(new_n760));
  INV_X1    g335(.A(G288), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n731), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT91), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT33), .B(G1976), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n731), .A2(G22), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G166), .B2(new_n731), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G1971), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(G1971), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n759), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT34), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT34), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n486), .A2(G119), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n481), .A2(G131), .ZN(new_n776));
  NOR2_X1   g351(.A1(G95), .A2(G2105), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(new_n477), .B2(G107), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G25), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT89), .B1(new_n781), .B2(G29), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n781), .A2(KEYINPUT89), .A3(G29), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT35), .B(G1991), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n731), .A2(G24), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G290), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1986), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n756), .B1(new_n774), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g370(.A(KEYINPUT36), .B(new_n793), .C1(new_n772), .C2(new_n773), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n750), .B(new_n755), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n587), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G4), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1348), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n731), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n540), .B2(new_n731), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G1341), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n797), .A2(new_n801), .A3(new_n805), .ZN(G311));
  NOR2_X1   g381(.A1(new_n795), .A2(new_n796), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n749), .ZN(new_n808));
  INV_X1    g383(.A(new_n801), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n808), .A2(new_n809), .A3(new_n804), .A4(new_n755), .ZN(G150));
  NAND2_X1  g385(.A1(new_n526), .A2(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n523), .A2(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n510), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n540), .B(new_n814), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n586), .A2(new_n594), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(G860), .ZN(G145));
  NAND3_X1  g397(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n491), .B1(new_n474), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n477), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n496), .A2(new_n497), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G2105), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n493), .A2(new_n494), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n713), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n745), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n832), .B2(new_n831), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n779), .B(new_n611), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n481), .A2(G142), .ZN(new_n837));
  NOR2_X1   g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G130), .B2(new_n486), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n835), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n607), .B(new_n479), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g424(.A(G303), .B(G288), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G305), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G290), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(KEYINPUT42), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT107), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(KEYINPUT42), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT106), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n596), .B(new_n817), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n587), .A2(new_n858), .A3(new_n736), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n736), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g435(.A1(G299), .A2(KEYINPUT105), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n586), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(KEYINPUT41), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(new_n857), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n854), .A2(new_n856), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n854), .B2(new_n856), .ZN(new_n870));
  OAI21_X1  g445(.A(G868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n814), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(G295));
  INV_X1    g449(.A(new_n870), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n872), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  INV_X1    g451(.A(new_n873), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT108), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n879), .A3(new_n873), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G331));
  XNOR2_X1  g456(.A(G168), .B(G301), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n817), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n863), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n865), .B2(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n885), .B2(new_n852), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n863), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n887), .B(new_n883), .C1(new_n865), .C2(KEYINPUT109), .ZN(new_n888));
  INV_X1    g463(.A(new_n884), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n886), .B1(new_n890), .B2(new_n852), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n885), .A2(new_n852), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT43), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT44), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n892), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(KEYINPUT43), .A3(new_n886), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n896), .B1(KEYINPUT44), .B2(new_n899), .ZN(G397));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(G164), .B2(G1384), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT110), .B(G40), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n472), .A2(new_n478), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G1996), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT111), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n909), .B(new_n911), .Z(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n745), .B(G2067), .Z(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n714), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(KEYINPUT127), .B2(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT47), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n713), .A2(G1996), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n913), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n714), .B2(new_n909), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n779), .A2(new_n786), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n745), .A2(G2067), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n906), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n779), .A2(new_n786), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n906), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(G290), .A2(new_n913), .A3(G1986), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT48), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n918), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G8), .ZN(new_n934));
  INV_X1    g509(.A(new_n905), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n829), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT115), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT50), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n937), .B2(KEYINPUT50), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n829), .A2(new_n944), .A3(new_n936), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n829), .B2(new_n936), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT114), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT113), .B1(G164), .B2(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n829), .A2(new_n944), .A3(new_n936), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n943), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n942), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n702), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n829), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n935), .B(new_n956), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n687), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n934), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G168), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT121), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT121), .B1(new_n959), .B2(G168), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n935), .B1(new_n945), .B2(new_n946), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(G1976), .B2(new_n761), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT119), .B(G1976), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n967), .B(new_n968), .C1(new_n761), .C2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(G305), .A2(G1981), .ZN(new_n971));
  NAND2_X1  g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(KEYINPUT49), .A3(new_n972), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979));
  INV_X1    g554(.A(G1976), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n980), .B2(G288), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n981), .B2(KEYINPUT52), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n967), .A2(KEYINPUT118), .A3(new_n968), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n970), .B(new_n978), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G166), .A2(new_n934), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT116), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT117), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT55), .B1(new_n986), .B2(KEYINPUT116), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n902), .A2(new_n956), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n935), .ZN(new_n993));
  INV_X1    g568(.A(G1971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n492), .A2(new_n498), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n996), .B2(new_n828), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT115), .B1(new_n997), .B2(new_n943), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n905), .B1(new_n998), .B2(new_n939), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n952), .B1(new_n951), .B2(new_n943), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n949), .C2(new_n950), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n995), .B1(new_n1002), .B2(G2090), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n991), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n990), .A2(G8), .A3(new_n1003), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n985), .A2(new_n1005), .A3(KEYINPUT63), .A4(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT63), .B1(new_n964), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1006), .A2(new_n984), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n978), .A2(new_n980), .A3(new_n761), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n976), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n955), .A2(G168), .A3(new_n958), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT51), .ZN(new_n1017));
  AOI21_X1  g592(.A(G168), .B1(new_n955), .B2(new_n958), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  OAI211_X1 g594(.A(G8), .B(new_n1015), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n954), .A2(G1961), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n993), .B2(G2078), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1022), .A2(G2078), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n957), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G301), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1017), .A2(new_n1020), .A3(KEYINPUT62), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n978), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT118), .B1(new_n967), .B2(new_n968), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n981), .A2(new_n979), .A3(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1006), .A2(new_n1032), .A3(KEYINPUT63), .A4(new_n970), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1005), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1028), .B1(new_n1035), .B2(new_n964), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1026), .A2(KEYINPUT62), .A3(G301), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n948), .A2(new_n953), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1348), .B1(new_n1039), .B2(new_n999), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n965), .A2(G2067), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n587), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(G299), .B(KEYINPUT57), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n949), .A2(KEYINPUT50), .A3(new_n950), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n905), .B1(new_n997), .B2(new_n943), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1956), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT56), .B(G2072), .ZN(new_n1047));
  AND4_X1   g622(.A1(new_n935), .A2(new_n902), .A3(new_n956), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1043), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1043), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(new_n1052), .C1(new_n1054), .C2(G1956), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1046), .A2(new_n1043), .A3(new_n1048), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT122), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1002), .A2(new_n800), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1041), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n586), .A2(KEYINPUT60), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n905), .B1(new_n949), .B2(new_n950), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT58), .B(G1341), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1068), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n965), .A2(KEYINPUT123), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n902), .A2(new_n935), .A3(new_n907), .A4(new_n956), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n540), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1073), .B2(new_n540), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1065), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1057), .A2(new_n1049), .A3(new_n1059), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1062), .A2(new_n586), .A3(new_n1063), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1042), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1058), .B1(KEYINPUT124), .B2(new_n1049), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n1046), .A2(new_n1048), .A3(new_n1043), .A4(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1084), .A2(new_n1078), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1061), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(G301), .B(KEYINPUT54), .Z(new_n1090));
  NOR3_X1   g665(.A1(new_n1021), .A2(new_n1025), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n954), .B2(G1961), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1002), .A2(KEYINPUT125), .A3(new_n722), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n992), .A2(G40), .A3(G160), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(new_n1024), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1093), .A2(new_n1023), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1091), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1038), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1036), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1053), .A2(KEYINPUT120), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n754), .B1(new_n1053), .B2(KEYINPUT120), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n995), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n985), .B(new_n1006), .C1(new_n990), .C2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1014), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(G290), .B(new_n790), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n928), .B1(new_n913), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1109), .B(KEYINPUT112), .Z(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT126), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n586), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n587), .B(new_n1041), .C1(new_n1002), .C2(new_n800), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1079), .A2(new_n1078), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1073), .A2(new_n540), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1073), .A2(new_n1074), .A3(new_n540), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1041), .B1(new_n1002), .B2(new_n800), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1117), .A2(new_n1118), .B1(new_n1119), .B2(new_n1064), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1055), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1086), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1114), .A2(new_n1115), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1098), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1100), .B1(new_n1127), .B2(new_n1037), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1017), .A2(new_n1020), .A3(KEYINPUT62), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n960), .B(new_n961), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1027), .B1(new_n1130), .B2(new_n1007), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1106), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT126), .B(new_n1110), .C1(new_n1132), .C2(new_n1013), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n933), .B1(new_n1111), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g710(.A(new_n899), .ZN(new_n1137));
  NOR3_X1   g711(.A1(G229), .A2(G401), .A3(G227), .ZN(new_n1138));
  NAND4_X1  g712(.A1(new_n1137), .A2(new_n1138), .A3(new_n462), .A4(new_n848), .ZN(G225));
  INV_X1    g713(.A(G225), .ZN(G308));
endmodule


