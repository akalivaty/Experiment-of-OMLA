

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579;

  XOR2_X1 U324 ( .A(n393), .B(n308), .Z(n545) );
  XOR2_X1 U325 ( .A(n425), .B(n424), .Z(n292) );
  XOR2_X1 U326 ( .A(G120GAT), .B(G127GAT), .Z(n293) );
  XOR2_X1 U327 ( .A(n306), .B(n305), .Z(n294) );
  NOR2_X1 U328 ( .A1(n555), .A2(n504), .ZN(n505) );
  INV_X1 U329 ( .A(KEYINPUT103), .ZN(n410) );
  XNOR2_X1 U330 ( .A(n426), .B(n292), .ZN(n427) );
  XNOR2_X1 U331 ( .A(n410), .B(KEYINPUT37), .ZN(n411) );
  XNOR2_X1 U332 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U333 ( .A(n412), .B(n411), .ZN(n487) );
  NOR2_X1 U334 ( .A1(n545), .A2(n544), .ZN(n556) );
  XNOR2_X1 U335 ( .A(KEYINPUT41), .B(n567), .ZN(n549) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n450) );
  XNOR2_X1 U337 ( .A(KEYINPUT38), .B(n449), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U340 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U342 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U344 ( .A(n297), .B(G183GAT), .Z(n299) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(G176GAT), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n393) );
  XNOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n293), .B(n300), .ZN(n359) );
  XOR2_X1 U349 ( .A(KEYINPUT20), .B(n359), .Z(n302) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U352 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U355 ( .A(G43GAT), .B(G15GAT), .Z(n432) );
  XOR2_X1 U356 ( .A(G99GAT), .B(G71GAT), .Z(n418) );
  XNOR2_X1 U357 ( .A(n432), .B(n418), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n294), .B(n307), .ZN(n308) );
  XOR2_X1 U359 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n318) );
  NAND2_X1 U362 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U363 ( .A(G211GAT), .B(G127GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(G22GAT), .B(G71GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n314) );
  XOR2_X1 U366 ( .A(G155GAT), .B(G78GAT), .Z(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n330) );
  XOR2_X1 U370 ( .A(G57GAT), .B(G183GAT), .Z(n320) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(G1GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(KEYINPUT13), .Z(n324) );
  XNOR2_X1 U377 ( .A(G8GAT), .B(G64GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U379 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n519) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G50GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n435) );
  XOR2_X1 U385 ( .A(G85GAT), .B(G92GAT), .Z(n416) );
  XOR2_X1 U386 ( .A(n435), .B(n416), .Z(n334) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U389 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT75), .B(KEYINPUT10), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U392 ( .A(n338), .B(n337), .Z(n346) );
  XOR2_X1 U393 ( .A(G218GAT), .B(G162GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(G134GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U396 ( .A(G106GAT), .B(G99GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n555) );
  XOR2_X1 U401 ( .A(n555), .B(KEYINPUT36), .Z(n577) );
  XNOR2_X1 U402 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n347), .B(KEYINPUT2), .ZN(n348) );
  XOR2_X1 U404 ( .A(n348), .B(KEYINPUT3), .Z(n350) );
  XNOR2_X1 U405 ( .A(G155GAT), .B(G162GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n383) );
  XOR2_X1 U407 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n352) );
  XNOR2_X1 U408 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n383), .B(n353), .ZN(n363) );
  XOR2_X1 U411 ( .A(G148GAT), .B(G57GAT), .Z(n415) );
  XOR2_X1 U412 ( .A(G1GAT), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U413 ( .A(G29GAT), .B(G141GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n431) );
  XOR2_X1 U415 ( .A(n415), .B(n431), .Z(n357) );
  NAND2_X1 U416 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n358), .B(KEYINPUT1), .Z(n361) );
  XNOR2_X1 U419 ( .A(n359), .B(KEYINPUT4), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n403) );
  XOR2_X1 U422 ( .A(G148GAT), .B(KEYINPUT22), .Z(n365) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U425 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n367) );
  XNOR2_X1 U426 ( .A(G22GAT), .B(G141GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U428 ( .A(n369), .B(n368), .Z(n381) );
  XNOR2_X1 U429 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n370), .B(KEYINPUT89), .ZN(n371) );
  XOR2_X1 U431 ( .A(n371), .B(KEYINPUT90), .Z(n373) );
  XNOR2_X1 U432 ( .A(G211GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n387) );
  XOR2_X1 U434 ( .A(G106GAT), .B(G78GAT), .Z(n417) );
  XOR2_X1 U435 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n375) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U438 ( .A(n417), .B(n376), .Z(n378) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n387), .B(n379), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n542) );
  XOR2_X1 U444 ( .A(G204GAT), .B(G64GAT), .Z(n413) );
  XOR2_X1 U445 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n385) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n413), .B(n386), .ZN(n391) );
  XOR2_X1 U449 ( .A(G92GAT), .B(n387), .Z(n389) );
  XOR2_X1 U450 ( .A(G197GAT), .B(G8GAT), .Z(n433) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(n433), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n538) );
  NOR2_X1 U455 ( .A1(n545), .A2(n538), .ZN(n394) );
  NOR2_X1 U456 ( .A1(n542), .A2(n394), .ZN(n395) );
  XOR2_X1 U457 ( .A(KEYINPUT25), .B(n395), .Z(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n396), .B(n538), .ZN(n404) );
  NAND2_X1 U460 ( .A1(n542), .A2(n545), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n397), .B(KEYINPUT100), .ZN(n398) );
  XNOR2_X1 U462 ( .A(KEYINPUT26), .B(n398), .ZN(n562) );
  NOR2_X1 U463 ( .A1(n404), .A2(n562), .ZN(n399) );
  NOR2_X1 U464 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U465 ( .A1(n403), .A2(n401), .ZN(n408) );
  XOR2_X1 U466 ( .A(n545), .B(KEYINPUT85), .Z(n402) );
  XOR2_X1 U467 ( .A(KEYINPUT28), .B(n542), .Z(n512) );
  NAND2_X1 U468 ( .A1(n402), .A2(n512), .ZN(n406) );
  XNOR2_X1 U469 ( .A(KEYINPUT95), .B(n403), .ZN(n540) );
  NOR2_X1 U470 ( .A1(n404), .A2(n540), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n405), .B(KEYINPUT99), .ZN(n511) );
  NOR2_X1 U472 ( .A1(n406), .A2(n511), .ZN(n407) );
  NOR2_X1 U473 ( .A1(n408), .A2(n407), .ZN(n454) );
  NOR2_X1 U474 ( .A1(n577), .A2(n454), .ZN(n409) );
  NAND2_X1 U475 ( .A1(n519), .A2(n409), .ZN(n412) );
  XNOR2_X1 U476 ( .A(G176GAT), .B(G120GAT), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n430) );
  XOR2_X1 U478 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n428) );
  XOR2_X1 U481 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n422) );
  XNOR2_X1 U482 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n423), .B(KEYINPUT72), .ZN(n426) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n425) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n567) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U490 ( .A(n435), .B(KEYINPUT69), .Z(n437) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(n439), .B(n438), .Z(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n441) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G22GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U497 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n443) );
  XNOR2_X1 U498 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n564) );
  XNOR2_X1 U502 ( .A(KEYINPUT70), .B(n564), .ZN(n546) );
  NAND2_X1 U503 ( .A1(n567), .A2(n546), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT74), .B(n448), .Z(n457) );
  NAND2_X1 U505 ( .A1(n487), .A2(n457), .ZN(n449) );
  NOR2_X1 U506 ( .A1(n545), .A2(n472), .ZN(n453) );
  XNOR2_X1 U507 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n451) );
  NOR2_X1 U508 ( .A1(n555), .A2(n519), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT16), .B(n455), .Z(n456) );
  NOR2_X1 U510 ( .A1(n454), .A2(n456), .ZN(n475) );
  NAND2_X1 U511 ( .A1(n475), .A2(n457), .ZN(n465) );
  NOR2_X1 U512 ( .A1(n540), .A2(n465), .ZN(n458) );
  XOR2_X1 U513 ( .A(G1GAT), .B(n458), .Z(n459) );
  XNOR2_X1 U514 ( .A(KEYINPUT34), .B(n459), .ZN(G1324GAT) );
  NOR2_X1 U515 ( .A1(n538), .A2(n465), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U518 ( .A(G8GAT), .B(n462), .ZN(G1325GAT) );
  NOR2_X1 U519 ( .A1(n545), .A2(n465), .ZN(n464) );
  XNOR2_X1 U520 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NOR2_X1 U522 ( .A1(n512), .A2(n465), .ZN(n466) );
  XOR2_X1 U523 ( .A(G22GAT), .B(n466), .Z(G1327GAT) );
  NOR2_X1 U524 ( .A1(n472), .A2(n540), .ZN(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(G29GAT), .B(n469), .ZN(G1328GAT) );
  NOR2_X1 U528 ( .A1(n472), .A2(n538), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(G1329GAT) );
  NOR2_X1 U531 ( .A1(n472), .A2(n512), .ZN(n473) );
  XOR2_X1 U532 ( .A(G50GAT), .B(n473), .Z(G1331GAT) );
  INV_X1 U533 ( .A(n549), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n564), .A2(n474), .ZN(n486) );
  NAND2_X1 U535 ( .A1(n486), .A2(n475), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT108), .B(n476), .ZN(n482) );
  NOR2_X1 U537 ( .A1(n482), .A2(n540), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G57GAT), .B(n479), .ZN(G1332GAT) );
  NOR2_X1 U541 ( .A1(n482), .A2(n538), .ZN(n480) );
  XOR2_X1 U542 ( .A(G64GAT), .B(n480), .Z(G1333GAT) );
  NOR2_X1 U543 ( .A1(n545), .A2(n482), .ZN(n481) );
  XOR2_X1 U544 ( .A(G71GAT), .B(n481), .Z(G1334GAT) );
  NOR2_X1 U545 ( .A1(n482), .A2(n512), .ZN(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U548 ( .A(G78GAT), .B(n485), .Z(G1335GAT) );
  NAND2_X1 U549 ( .A1(n487), .A2(n486), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n540), .A2(n492), .ZN(n488) );
  XOR2_X1 U551 ( .A(G85GAT), .B(n488), .Z(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT110), .B(n489), .ZN(G1336GAT) );
  NOR2_X1 U553 ( .A1(n538), .A2(n492), .ZN(n490) );
  XOR2_X1 U554 ( .A(G92GAT), .B(n490), .Z(G1337GAT) );
  NOR2_X1 U555 ( .A1(n545), .A2(n492), .ZN(n491) );
  XOR2_X1 U556 ( .A(G99GAT), .B(n491), .Z(G1338GAT) );
  NOR2_X1 U557 ( .A1(n512), .A2(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n495), .ZN(G1339GAT) );
  XNOR2_X1 U561 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n516) );
  XOR2_X1 U562 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n497) );
  NOR2_X1 U563 ( .A1(n519), .A2(n577), .ZN(n496) );
  XOR2_X1 U564 ( .A(n497), .B(n496), .Z(n498) );
  NAND2_X1 U565 ( .A1(n567), .A2(n498), .ZN(n499) );
  NOR2_X1 U566 ( .A1(n546), .A2(n499), .ZN(n500) );
  XOR2_X1 U567 ( .A(KEYINPUT115), .B(n500), .Z(n509) );
  XOR2_X1 U568 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n501) );
  XNOR2_X1 U569 ( .A(KEYINPUT112), .B(n501), .ZN(n503) );
  NAND2_X1 U570 ( .A1(n549), .A2(n564), .ZN(n502) );
  XOR2_X1 U571 ( .A(n503), .B(n502), .Z(n504) );
  NAND2_X1 U572 ( .A1(n505), .A2(n519), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(KEYINPUT114), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT47), .ZN(n508) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT48), .B(n510), .ZN(n537) );
  OR2_X1 U577 ( .A1(n537), .A2(n511), .ZN(n525) );
  INV_X1 U578 ( .A(n545), .ZN(n513) );
  NAND2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n514) );
  NOR2_X1 U580 ( .A1(n525), .A2(n514), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n546), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U584 ( .A1(n522), .A2(n549), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  INV_X1 U586 ( .A(n519), .ZN(n572) );
  NAND2_X1 U587 ( .A1(n572), .A2(n522), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(KEYINPUT50), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(n521), .ZN(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n555), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  XNOR2_X1 U593 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n562), .A2(n525), .ZN(n526) );
  XOR2_X1 U595 ( .A(KEYINPUT117), .B(n526), .Z(n535) );
  NAND2_X1 U596 ( .A1(n564), .A2(n535), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(G1344GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n530) );
  NAND2_X1 U599 ( .A1(n535), .A2(n549), .ZN(n529) );
  XNOR2_X1 U600 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT53), .Z(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(G1345GAT) );
  NAND2_X1 U603 ( .A1(n572), .A2(n535), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n533), .B(KEYINPUT120), .ZN(n534) );
  XNOR2_X1 U605 ( .A(G155GAT), .B(n534), .ZN(G1346GAT) );
  NAND2_X1 U606 ( .A1(n535), .A2(n555), .ZN(n536) );
  XNOR2_X1 U607 ( .A(n536), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U608 ( .A(G169GAT), .B(KEYINPUT121), .Z(n548) );
  NOR2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n539), .B(KEYINPUT54), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n563) );
  NOR2_X1 U612 ( .A1(n563), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n543), .B(KEYINPUT55), .ZN(n544) );
  NAND2_X1 U614 ( .A1(n556), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1348GAT) );
  XNOR2_X1 U616 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n556), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n550) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1349GAT) );
  NAND2_X1 U620 ( .A1(n572), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT58), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(n558), .ZN(G1351GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n560) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(n561), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n573), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  INV_X1 U632 ( .A(n573), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n576), .A2(n567), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n569) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  XOR2_X1 U638 ( .A(G211GAT), .B(KEYINPUT127), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

