//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT66), .Z(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT67), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n222), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n207), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n219), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT74), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G20), .A2(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT15), .B(G87), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n228), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n251), .B1(new_n252), .B2(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n227), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n264), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n259), .B1(new_n263), .B2(new_n265), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(G77), .C1(G1), .C2(new_n228), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n260), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(KEYINPUT69), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G232), .ZN(new_n281));
  INV_X1    g0081(.A(G238), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n281), .C1(new_n282), .C2(new_n280), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n278), .B(new_n283), .C1(G107), .C2(new_n279), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n276), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(G244), .ZN(new_n291));
  AOI21_X1  g0091(.A(G169), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n250), .B1(new_n271), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n284), .A2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n260), .A2(new_n268), .A3(new_n270), .ZN(new_n297));
  OAI211_X1 g0097(.A(KEYINPUT74), .B(new_n297), .C1(new_n294), .C2(G169), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(G58), .B(G68), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT7), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n279), .B2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT7), .B(new_n228), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT77), .B1(new_n310), .B2(G68), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT77), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n304), .C2(new_n309), .ZN(new_n314));
  OAI211_X1 g0114(.A(KEYINPUT16), .B(new_n302), .C1(new_n311), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(G68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n302), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n259), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n269), .B1(G1), .B2(new_n228), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT70), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n256), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n266), .B2(new_n324), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n327));
  OR2_X1    g0127(.A1(G223), .A2(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n305), .A2(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n217), .A2(G1698), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n287), .B1(new_n278), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n290), .A2(G232), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n334), .A2(new_n336), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n321), .A2(new_n326), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n321), .A2(new_n326), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n321), .A2(new_n326), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n334), .A2(G179), .A3(new_n336), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n334), .B2(new_n336), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT18), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n352), .B(new_n349), .C1(new_n321), .C2(new_n326), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n341), .A2(new_n344), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT80), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n300), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n327), .A2(new_n329), .A3(G232), .A4(G1698), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n279), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n360));
  AND2_X1   g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n360), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n278), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n285), .A2(new_n286), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n289), .B2(new_n282), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT13), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(G190), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n365), .B2(new_n368), .ZN(new_n374));
  AOI211_X1 g0174(.A(KEYINPUT13), .B(new_n367), .C1(new_n364), .C2(new_n278), .ZN(new_n375));
  OAI21_X1  g0175(.A(G200), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n307), .A2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G77), .B1(G20), .B2(new_n313), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n216), .B2(new_n255), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n259), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT11), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT11), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n382), .A3(new_n259), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n263), .A2(new_n265), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n322), .A2(new_n313), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n373), .A2(new_n376), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT76), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n373), .A2(new_n376), .A3(new_n391), .A4(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n374), .B2(new_n375), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n374), .A2(new_n375), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(G169), .C1(new_n374), .C2(new_n375), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n390), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n294), .A2(new_n405), .ZN(new_n406));
  OR3_X1    g0206(.A1(new_n297), .A2(new_n406), .A3(KEYINPUT73), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n294), .A2(G190), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT73), .B1(new_n406), .B2(new_n297), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n396), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n353), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n345), .A2(new_n350), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n352), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n343), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(KEYINPUT80), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n280), .A2(G222), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G223), .A2(G1698), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n279), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n278), .B(new_n421), .C1(G77), .C2(new_n279), .ZN(new_n422));
  OR2_X1    g0222(.A1(KEYINPUT68), .A2(G226), .ZN(new_n423));
  NAND2_X1  g0223(.A1(KEYINPUT68), .A2(G226), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n290), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n366), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n216), .B1(new_n261), .B2(G20), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n428), .A2(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(KEYINPUT72), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n269), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n432));
  INV_X1    g0232(.A(G150), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n255), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n324), .B2(new_n377), .ZN(new_n435));
  INV_X1    g0235(.A(new_n259), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n431), .B1(G50), .B2(new_n385), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n347), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n427), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n426), .A2(G200), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n440), .B1(new_n335), .B2(new_n426), .C1(new_n437), .C2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n437), .A2(new_n441), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT10), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT10), .B1(new_n442), .B2(new_n443), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n356), .A2(new_n411), .A3(new_n418), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n261), .A2(G33), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n269), .A2(G116), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n266), .A2(new_n218), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n258), .A2(new_n227), .B1(G20), .B2(new_n218), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n228), .C1(G33), .C2(new_n212), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT20), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n453), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n449), .B(new_n450), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n327), .A2(new_n329), .ZN(new_n457));
  INV_X1    g0257(.A(G303), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G264), .A2(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n279), .B(new_n460), .C1(new_n213), .C2(G1698), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n278), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n261), .B(G45), .C1(new_n463), .C2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT83), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n261), .A4(G45), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(G274), .C1(new_n273), .C2(new_n227), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n466), .A2(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n288), .B(G270), .C1(new_n464), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n462), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n456), .A2(new_n477), .A3(G169), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT21), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n456), .A2(new_n477), .A3(new_n480), .A4(G169), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT87), .ZN(new_n482));
  INV_X1    g0282(.A(new_n456), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n462), .A2(G179), .A3(new_n474), .A4(new_n476), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n484), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT87), .A3(new_n456), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n479), .A2(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n327), .A2(new_n329), .A3(new_n228), .A4(G87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n279), .A2(new_n228), .A3(G87), .A4(new_n490), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n228), .A2(G107), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT23), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n494), .A2(KEYINPUT24), .A3(new_n495), .A4(new_n497), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n259), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n269), .A2(new_n448), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n385), .A2(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT25), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT89), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n274), .A2(new_n277), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n211), .A2(new_n280), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n213), .A2(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n327), .A2(new_n511), .A3(new_n329), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n288), .B(G264), .C1(new_n464), .C2(new_n475), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n508), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n510), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n278), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n515), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n520), .A3(G179), .A4(new_n474), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n474), .A3(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n507), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n477), .A2(G200), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n483), .C1(new_n335), .C2(new_n477), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n488), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(new_n520), .A3(new_n474), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n405), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n522), .A2(G190), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n261), .A2(G45), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n211), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n288), .C1(G274), .C2(new_n535), .ZN(new_n537));
  MUX2_X1   g0337(.A(G238), .B(G244), .S(G1698), .Z(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n279), .B1(G33), .B2(G116), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n509), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n295), .ZN(new_n542));
  INV_X1    g0342(.A(new_n252), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n269), .A2(new_n543), .A3(new_n448), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n266), .A2(new_n252), .ZN(new_n545));
  NOR3_X1   g0345(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n361), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n546), .B1(new_n551), .B2(new_n228), .ZN(new_n552));
  AOI22_X1  g0352(.A1(G97), .A2(new_n377), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  AND4_X1   g0353(.A1(new_n228), .A2(new_n327), .A3(new_n329), .A4(G68), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n544), .B(new_n545), .C1(new_n555), .C2(new_n436), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n540), .A2(new_n347), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n542), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n269), .A2(G87), .A3(new_n448), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n269), .A2(KEYINPUT86), .A3(G87), .A4(new_n448), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n253), .A2(new_n212), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n279), .A2(new_n228), .A3(G68), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n564), .A2(new_n565), .ZN(new_n568));
  AOI21_X1  g0368(.A(G20), .B1(new_n568), .B2(new_n361), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n567), .C1(new_n569), .C2(new_n546), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n259), .B1(new_n266), .B2(new_n252), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n540), .A2(G200), .ZN(new_n572));
  OAI211_X1 g0372(.A(G190), .B(new_n537), .C1(new_n539), .C2(new_n509), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n563), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n558), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n385), .B2(G97), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n212), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(new_n503), .B2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT7), .B1(new_n457), .B2(new_n228), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n303), .B(G20), .C1(new_n327), .C2(new_n329), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  AND2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G97), .A2(G107), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(KEYINPUT6), .A3(G97), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n580), .B1(new_n592), .B2(new_n259), .ZN(new_n593));
  AOI211_X1 g0393(.A(KEYINPUT81), .B(new_n436), .C1(new_n583), .C2(new_n591), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n579), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n327), .A2(new_n329), .A3(G244), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n599), .A3(new_n452), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n279), .A2(G250), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n280), .B1(new_n601), .B2(KEYINPUT4), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n278), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n472), .B1(new_n469), .B2(new_n465), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n288), .B(G257), .C1(new_n464), .C2(new_n475), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n606), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n347), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n295), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n595), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n589), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n584), .B2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n228), .B1(new_n267), .B2(new_n255), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n588), .B1(new_n304), .B2(new_n309), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n259), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n592), .A2(new_n580), .A3(new_n259), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n610), .A2(G200), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n603), .A2(new_n608), .A3(new_n609), .A4(G190), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n579), .A4(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n534), .A2(new_n575), .A3(new_n614), .A4(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n447), .A2(new_n528), .A3(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n444), .A2(new_n445), .ZN(new_n629));
  INV_X1    g0429(.A(new_n417), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n390), .B1(new_n399), .B2(G190), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT76), .B1(new_n631), .B2(new_n376), .ZN(new_n632));
  INV_X1    g0432(.A(new_n395), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n300), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n634), .B2(new_n404), .ZN(new_n635));
  INV_X1    g0435(.A(new_n415), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n439), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n447), .ZN(new_n640));
  INV_X1    g0440(.A(new_n558), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n558), .A2(new_n574), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n614), .B2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n623), .A2(new_n579), .B1(new_n347), .B2(new_n610), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n575), .A3(KEYINPUT26), .A4(new_n613), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n641), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n525), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n507), .A2(KEYINPUT90), .A3(new_n524), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n649), .A2(new_n488), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n627), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n639), .B1(new_n640), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT91), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n261), .A2(new_n228), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(KEYINPUT92), .A2(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(KEYINPUT92), .A2(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n483), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n488), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n488), .A2(new_n527), .A3(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT93), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n507), .A2(new_n524), .A3(new_n663), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT95), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT94), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n529), .B2(new_n664), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n507), .A2(KEYINPUT94), .A3(new_n663), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n525), .A3(new_n534), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT96), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n674), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n672), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n488), .A2(new_n663), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n680), .B2(new_n682), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n663), .B1(new_n649), .B2(new_n650), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n204), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n546), .A2(new_n218), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n232), .B2(new_n695), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n517), .A2(new_n520), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n612), .A3(new_n486), .A4(new_n541), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n610), .A2(new_n295), .A3(new_n477), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n530), .A3(new_n540), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n663), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n627), .A2(new_n528), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n664), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n663), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n534), .A2(new_n614), .A3(new_n626), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n649), .A2(new_n488), .A3(new_n650), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n575), .ZN(new_n719));
  AOI211_X1 g0519(.A(KEYINPUT29), .B(new_n663), .C1(new_n719), .C2(new_n647), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n614), .A2(new_n626), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n488), .A2(new_n525), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n723), .A3(new_n575), .A4(new_n534), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n647), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n725), .B2(new_n664), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n716), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n700), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n695), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n672), .B(new_n734), .C1(G330), .C2(new_n669), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n227), .B1(G20), .B2(new_n347), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n228), .A2(new_n295), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(G190), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n228), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n335), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G326), .A2(new_n740), .B1(new_n743), .B2(G283), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n228), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G329), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n744), .B(new_n749), .C1(new_n458), .C2(new_n750), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n228), .A2(new_n295), .A3(G190), .A4(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n738), .A2(new_n335), .A3(G200), .ZN(new_n756));
  OR2_X1    g0556(.A1(KEYINPUT33), .A2(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(KEYINPUT33), .A2(G317), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n751), .A2(new_n279), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n228), .B1(new_n746), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n738), .A2(G190), .A3(new_n405), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT100), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT100), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n738), .A2(new_n766), .A3(G190), .A4(new_n405), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n763), .C2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT101), .Z(new_n771));
  NAND2_X1  g0571(.A1(new_n748), .A2(G159), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n279), .B1(new_n739), .B2(new_n216), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n750), .A2(new_n210), .ZN(new_n776));
  INV_X1    g0576(.A(G58), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n753), .A2(new_n267), .B1(new_n762), .B2(new_n212), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n780), .B1(new_n313), .B2(new_n756), .C1(new_n588), .C2(new_n742), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n737), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n736), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT99), .Z(new_n787));
  NAND3_X1  g0587(.A1(new_n279), .A2(G355), .A3(new_n204), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G116), .B2(new_n204), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  INV_X1    g0590(.A(G45), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n233), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n693), .A2(new_n279), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(new_n245), .C2(new_n791), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n787), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n782), .A2(new_n795), .A3(new_n734), .ZN(new_n796));
  INV_X1    g0596(.A(new_n785), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n669), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n735), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  OAI22_X1  g0600(.A1(new_n753), .A2(new_n218), .B1(new_n458), .B2(new_n739), .ZN(new_n801));
  INV_X1    g0601(.A(new_n756), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G283), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT102), .Z(new_n804));
  AOI211_X1 g0604(.A(new_n279), .B(new_n804), .C1(G311), .C2(new_n748), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n805), .B1(new_n210), .B2(new_n742), .C1(new_n588), .C2(new_n750), .ZN(new_n806));
  INV_X1    g0606(.A(new_n762), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n768), .A2(G294), .B1(G97), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT103), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n279), .B1(new_n762), .B2(new_n777), .C1(new_n810), .C2(new_n747), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n768), .A2(G143), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n740), .B1(new_n802), .B2(G150), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n753), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n816), .B1(new_n216), .B2(new_n750), .C1(new_n313), .C2(new_n742), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n806), .A2(new_n809), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n736), .A2(new_n783), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(new_n736), .B1(new_n267), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n299), .A2(KEYINPUT104), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT104), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n293), .A2(new_n298), .A3(new_n822), .A4(new_n296), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n297), .A2(new_n663), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n824), .A2(new_n410), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n299), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n784), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n734), .B1(new_n820), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n652), .A2(new_n664), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(new_n828), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(new_n716), .ZN(new_n835));
  INV_X1    g0635(.A(new_n734), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT105), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT108), .ZN(new_n840));
  INV_X1    g0640(.A(new_n658), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n345), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n413), .A2(new_n842), .A3(new_n844), .A4(new_n340), .ZN(new_n845));
  INV_X1    g0645(.A(new_n340), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n321), .A2(new_n326), .B1(new_n349), .B2(new_n658), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n354), .A2(new_n843), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n849), .B2(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(new_n302), .ZN(new_n851));
  INV_X1    g0651(.A(new_n311), .ZN(new_n852));
  INV_X1    g0652(.A(new_n314), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n259), .B(new_n315), .C1(new_n854), .C2(new_n318), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(new_n326), .B1(new_n349), .B2(new_n658), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n856), .B2(new_n846), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n845), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT107), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n326), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n354), .A2(new_n841), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(new_n845), .A3(KEYINPUT107), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT38), .A4(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n842), .B1(new_n415), .B2(new_n417), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n845), .A2(new_n848), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT108), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n850), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n488), .A2(new_n525), .A3(new_n527), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n717), .A2(new_n870), .A3(new_n575), .A4(new_n664), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n396), .A2(new_n404), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n390), .A2(new_n663), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n396), .A2(new_n404), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n872), .A2(new_n878), .A3(new_n710), .A4(new_n828), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n879), .A3(KEYINPUT40), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n865), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n864), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT40), .B1(new_n884), .B2(new_n879), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n640), .A2(new_n715), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G330), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n652), .A2(new_n664), .A3(new_n828), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n824), .A2(new_n663), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n895), .A2(new_n884), .B1(new_n636), .B2(new_n658), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n869), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n404), .A2(new_n663), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n864), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n889), .B(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n652), .A2(new_n721), .A3(new_n664), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n663), .B1(new_n724), .B2(new_n647), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n721), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n639), .B1(new_n906), .B2(new_n640), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n903), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n261), .B2(new_n732), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n218), .B1(new_n590), .B2(KEYINPUT35), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n910), .B(new_n229), .C1(KEYINPUT35), .C2(new_n590), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n777), .B2(new_n313), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n232), .A2(new_n913), .B1(G50), .B2(new_n313), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n731), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(G367));
  AOI21_X1  g0716(.A(new_n279), .B1(new_n748), .B2(G317), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n743), .A2(G97), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n918), .C1(new_n754), .C2(new_n739), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G107), .B2(new_n807), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n768), .A2(G303), .ZN(new_n921));
  INV_X1    g0721(.A(new_n750), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G116), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n802), .A2(G294), .B1(G283), .B2(new_n752), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n920), .A2(new_n921), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G143), .A2(new_n740), .B1(new_n922), .B2(G58), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n216), .B2(new_n753), .C1(new_n313), .C2(new_n762), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n457), .B(new_n928), .C1(G159), .C2(new_n802), .ZN(new_n929));
  INV_X1    g0729(.A(G137), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n929), .B1(new_n267), .B2(new_n742), .C1(new_n930), .C2(new_n747), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n769), .A2(new_n433), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n736), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n664), .B1(new_n563), .B2(new_n571), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n641), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n643), .B2(new_n936), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(new_n797), .ZN(new_n939));
  INV_X1    g0739(.A(new_n793), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n786), .B1(new_n204), .B2(new_n252), .C1(new_n241), .C2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n935), .A2(new_n836), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n733), .A2(G1), .ZN(new_n943));
  INV_X1    g0743(.A(new_n595), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n722), .B1(new_n944), .B2(new_n664), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n645), .A2(new_n613), .A3(new_n663), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT45), .B1(new_n691), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  INV_X1    g0749(.A(new_n947), .ZN(new_n950));
  NOR4_X1   g0750(.A1(new_n689), .A2(new_n949), .A3(new_n690), .A4(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT44), .B1(new_n691), .B2(new_n947), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n953), .A2(new_n686), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n685), .B1(new_n957), .B2(new_n952), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n683), .A2(new_n687), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n689), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n671), .A2(KEYINPUT112), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n960), .B(new_n961), .Z(new_n962));
  NAND4_X1  g0762(.A1(new_n956), .A2(new_n958), .A3(new_n729), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n729), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n694), .B(KEYINPUT41), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n943), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n689), .A2(new_n947), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n614), .B1(new_n945), .B2(new_n525), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n664), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT109), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT110), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n976), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n977), .A2(new_n976), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n972), .A2(new_n979), .A3(new_n980), .A4(new_n974), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT111), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n685), .A2(new_n947), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n978), .B(new_n981), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n978), .A2(new_n982), .A3(new_n981), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n942), .B1(new_n966), .B2(new_n988), .ZN(G387));
  NAND3_X1  g0789(.A1(new_n696), .A2(new_n204), .A3(new_n279), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n238), .A2(new_n791), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n256), .A2(G50), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n992), .B(new_n993), .Z(new_n994));
  NAND2_X1  g0794(.A1(G68), .A2(G77), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n697), .A2(new_n791), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n793), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n990), .B1(G107), .B2(new_n204), .C1(new_n991), .C2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n753), .A2(new_n313), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n324), .A2(new_n802), .B1(G159), .B2(new_n740), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n807), .A2(new_n543), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n216), .C2(new_n769), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(G150), .C2(new_n748), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n922), .A2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1004), .A2(new_n279), .A3(new_n918), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n768), .A2(G317), .B1(G303), .B2(new_n752), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n754), .B2(new_n756), .C1(new_n763), .C2(new_n739), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT48), .ZN(new_n1009));
  INV_X1    g0809(.A(G283), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n762), .C1(new_n761), .C2(new_n750), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n279), .B1(new_n748), .B2(G326), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n218), .B2(new_n742), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1006), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT115), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n836), .B1(new_n787), .B2(new_n999), .C1(new_n1017), .C2(new_n737), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n684), .B2(new_n785), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n943), .B2(new_n962), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n962), .A2(new_n729), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n962), .A2(new_n729), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n694), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(G393));
  NAND2_X1  g0824(.A1(new_n956), .A2(new_n958), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1022), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n694), .A3(new_n963), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n956), .A2(new_n958), .A3(new_n943), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n768), .A2(G311), .B1(G317), .B2(new_n740), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT52), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n279), .B(new_n1030), .C1(G283), .C2(new_n922), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n761), .B2(new_n753), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n747), .A2(new_n763), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n762), .A2(new_n218), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n756), .A2(new_n458), .B1(new_n742), .B2(new_n588), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n753), .A2(new_n256), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n768), .A2(G159), .B1(G150), .B2(new_n740), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT51), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n748), .A2(G143), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n762), .A2(new_n267), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n457), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G50), .A2(new_n802), .B1(new_n743), .B2(G87), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1037), .B(new_n1044), .C1(G68), .C2(new_n922), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n736), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n950), .A2(new_n785), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n786), .B1(new_n212), .B2(new_n204), .C1(new_n248), .C2(new_n940), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n836), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1028), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1027), .A2(new_n1050), .ZN(G390));
  INV_X1    g0851(.A(new_n869), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n891), .B1(new_n905), .B2(new_n828), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n878), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1053), .A2(new_n1054), .B1(new_n404), .B2(new_n663), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n715), .A2(G330), .A3(new_n828), .A4(new_n878), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n898), .A2(new_n900), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n899), .B1(new_n894), .B2(new_n878), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1056), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1057), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n898), .B2(new_n900), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n943), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1058), .A2(new_n784), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n324), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n819), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n753), .A2(new_n212), .B1(new_n313), .B2(new_n742), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1041), .B(new_n1070), .C1(G283), .C2(new_n740), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n802), .A2(G107), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n768), .A2(G116), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n279), .B(new_n776), .C1(G294), .C2(new_n748), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT54), .B(G143), .Z(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n753), .A2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n279), .B1(new_n742), .B2(new_n216), .C1(new_n930), .C2(new_n756), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G159), .C2(new_n807), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n740), .A2(G128), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n748), .A2(G125), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n768), .A2(G132), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n922), .A2(G150), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT53), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1075), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n736), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1067), .A2(new_n836), .A3(new_n1069), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n396), .A2(new_n300), .B1(new_n390), .B2(new_n403), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n415), .B1(new_n1091), .B2(new_n630), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n439), .B1(new_n1092), .B2(new_n629), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n727), .B2(new_n447), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n872), .A2(new_n710), .ZN(new_n1095));
  INV_X1    g0895(.A(G330), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(new_n447), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT116), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT116), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n640), .A2(G330), .A3(new_n715), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n907), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n872), .A2(new_n710), .A3(G330), .A4(new_n828), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1054), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1057), .A2(new_n1104), .A3(new_n1053), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n894), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1057), .B2(new_n1104), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1065), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n695), .B1(new_n1065), .B2(new_n1109), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1090), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G378));
  NAND4_X1  g0913(.A1(new_n872), .A2(new_n878), .A3(new_n710), .A4(new_n828), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n864), .B2(new_n883), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n880), .B(G330), .C1(new_n1115), .C2(KEYINPUT40), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n901), .A3(new_n896), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n901), .B2(new_n896), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n446), .B(KEYINPUT119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n437), .A2(new_n841), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1118), .A2(new_n1119), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n902), .A2(new_n886), .A3(G330), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1130), .B2(new_n1117), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n943), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n734), .B1(new_n1127), .B2(new_n783), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(G33), .A2(G41), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT117), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n216), .C1(G41), .C2(new_n279), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n753), .A2(new_n930), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1077), .A2(new_n750), .B1(new_n1138), .B2(new_n739), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(G128), .C2(new_n768), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n810), .B2(new_n756), .C1(new_n433), .C2(new_n762), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT59), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1135), .B1(G124), .B2(new_n748), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n814), .B2(new_n742), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n769), .A2(new_n588), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1005), .B1(new_n218), .B2(new_n739), .C1(new_n252), .C2(new_n753), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n756), .A2(new_n212), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n742), .A2(new_n777), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G41), .B(new_n279), .C1(new_n807), .C2(G68), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n1010), .C2(new_n747), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n736), .B1(new_n1145), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n819), .A2(new_n216), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1133), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1132), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1060), .A2(new_n1159), .A3(new_n1064), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(KEYINPUT57), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n694), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1128), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1130), .A2(new_n1117), .A3(new_n1127), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(new_n1161), .B2(new_n1159), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT57), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1158), .B1(new_n1164), .B2(new_n1168), .ZN(G375));
  NAND2_X1  g0969(.A1(new_n1160), .A2(new_n943), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1054), .A2(new_n783), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n819), .A2(new_n313), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n753), .A2(new_n588), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1002), .B1(new_n761), .B2(new_n739), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G116), .C2(new_n802), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n457), .B1(new_n750), .B2(new_n212), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G77), .B2(new_n743), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n1010), .C2(new_n769), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G303), .B2(new_n748), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n753), .A2(new_n433), .B1(new_n777), .B2(new_n742), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n457), .B(new_n1180), .C1(G128), .C2(new_n748), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n739), .A2(new_n810), .B1(new_n762), .B2(new_n216), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n768), .B2(G137), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n756), .C2(new_n1077), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G159), .B2(new_n922), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n736), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1171), .A2(new_n836), .A3(new_n1172), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1170), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n965), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1109), .B2(new_n1191), .ZN(G381));
  NAND2_X1  g0992(.A1(new_n1132), .A2(new_n1157), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n695), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1162), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n838), .A3(new_n1112), .ZN(new_n1199));
  OR3_X1    g0999(.A1(G390), .A2(G393), .A3(G396), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1199), .A2(G387), .A3(new_n1200), .A4(G381), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT120), .Z(G407));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1112), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G407), .B(G213), .C1(new_n661), .C2(new_n1203), .ZN(G409));
  INV_X1    g1004(.A(KEYINPUT126), .ZN(new_n1205));
  INV_X1    g1005(.A(G390), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(G387), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G390), .B(new_n942), .C1(new_n966), .C2(new_n988), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(G387), .A2(KEYINPUT124), .A3(new_n1206), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(G393), .B(G396), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1207), .A2(new_n1212), .A3(new_n1208), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT125), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT125), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1207), .A2(new_n1212), .A3(new_n1208), .A4(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n662), .A2(G213), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(G2897), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1190), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1108), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n694), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT121), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(KEYINPUT121), .A3(new_n694), .A4(new_n1225), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1230), .B2(new_n1189), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n838), .B(new_n1188), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1221), .A2(KEYINPUT123), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1222), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1222), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1234), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1231), .A2(new_n1232), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1167), .A2(new_n965), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1158), .A2(new_n1112), .A3(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1220), .B(new_n1241), .C1(new_n1198), .C2(new_n1112), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1230), .A2(new_n1189), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n838), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1230), .A2(G384), .A3(new_n1189), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT62), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1221), .B1(G375), .B2(G378), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT62), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1233), .A4(new_n1241), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1219), .B1(new_n1243), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1242), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1245), .A2(new_n1234), .A3(new_n1246), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1236), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(KEYINPUT122), .A3(new_n1220), .A4(new_n1241), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1233), .A2(new_n1222), .A3(new_n1234), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1256), .A2(new_n1258), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT63), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1249), .A2(new_n1264), .A3(new_n1233), .A4(new_n1241), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  AND4_X1   g1066(.A1(new_n1254), .A2(new_n1262), .A3(new_n1266), .A4(new_n1219), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1205), .B1(new_n1253), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1258), .A2(new_n1261), .A3(new_n1242), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(new_n1254), .A3(new_n1248), .A4(new_n1251), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(new_n1214), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1262), .A2(new_n1266), .A3(new_n1219), .A4(new_n1254), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1268), .A2(new_n1273), .ZN(G405));
  NOR2_X1   g1074(.A1(new_n1219), .A2(KEYINPUT127), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1259), .A2(new_n1203), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1233), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1219), .A2(KEYINPUT127), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(G402));
endmodule


