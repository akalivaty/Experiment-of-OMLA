//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G469), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT3), .A4(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n204), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n203), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n204), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n219), .B2(new_n205), .ZN(new_n220));
  INV_X1    g034(.A(new_n210), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n206), .A2(G104), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n209), .B2(new_n210), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n222), .B(KEYINPUT4), .C1(new_n224), .C2(new_n204), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n197), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n195), .A2(G143), .ZN(new_n228));
  OAI211_X1 g042(.A(G128), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n196), .B(new_n198), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n217), .B1(new_n209), .B2(new_n210), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n219), .B2(new_n223), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n216), .A2(new_n225), .B1(new_n236), .B2(KEYINPUT10), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n242), .A3(new_n246), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n222), .A2(new_n231), .A3(new_n229), .A4(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n250), .B2(new_n253), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n237), .B(new_n249), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT80), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT80), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n249), .A4(new_n237), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n248), .A2(KEYINPUT81), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n222), .A2(new_n234), .B1(new_n231), .B2(new_n229), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n236), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT12), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n264), .B(new_n268), .C1(new_n236), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n194), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n194), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT82), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n249), .B1(new_n260), .B2(new_n237), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n193), .B1(new_n258), .B2(new_n262), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n189), .B(new_n272), .C1(new_n274), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n194), .B1(new_n263), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n270), .B(new_n193), .C1(new_n258), .C2(new_n262), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n189), .B(new_n280), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n189), .A2(new_n280), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G122), .ZN(new_n293));
  INV_X1    g107(.A(G113), .ZN(new_n294));
  INV_X1    g108(.A(G116), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G119), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(G119), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n294), .A2(KEYINPUT2), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G113), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n298), .A2(new_n302), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n222), .A3(new_n234), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT84), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n233), .A2(new_n235), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n308), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n307), .A2(new_n303), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n303), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n211), .A2(new_n213), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n215), .A3(G101), .ZN(new_n320));
  AND4_X1   g134(.A1(new_n315), .A2(new_n225), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n214), .A2(new_n215), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n322), .B2(new_n225), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n293), .B(new_n314), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n293), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n309), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n311), .A2(new_n308), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n229), .A2(new_n330), .A3(new_n231), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n330), .B2(new_n203), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT7), .B1(new_n333), .B2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n336), .C1(new_n330), .C2(new_n203), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT88), .B1(new_n340), .B2(new_n280), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n342), .B(G902), .C1(new_n324), .C2(new_n339), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n333), .A2(G953), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT86), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n332), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT6), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n314), .B1(new_n321), .B2(new_n323), .ZN(new_n352));
  INV_X1    g166(.A(new_n293), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n350), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n292), .B1(new_n344), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n310), .A2(new_n313), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n225), .A2(new_n318), .A3(new_n320), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT83), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n322), .A2(new_n315), .A3(new_n225), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n349), .B1(new_n363), .B2(new_n293), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n293), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n356), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n347), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n329), .A2(new_n338), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n363), .B2(new_n293), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n342), .B1(new_n370), .B2(G902), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n340), .A2(KEYINPUT88), .A3(new_n280), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n291), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n290), .B1(new_n358), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G113), .B(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT91), .B(G104), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(KEYINPUT65), .A2(G237), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT65), .A2(G237), .ZN(new_n381));
  AOI21_X1  g195(.A(G953), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n197), .A2(KEYINPUT89), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G143), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(G214), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT65), .A2(G237), .ZN(new_n388));
  NOR2_X1   g202(.A1(KEYINPUT65), .A2(G237), .ZN(new_n389));
  OAI211_X1 g203(.A(G214), .B(new_n191), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n385), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n246), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT17), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n391), .A3(new_n246), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G140), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n330), .B2(KEYINPUT72), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G125), .A3(G140), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(G125), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n401), .A2(new_n195), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n195), .B1(new_n401), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n392), .A2(KEYINPUT17), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n387), .A2(new_n391), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT18), .A3(G131), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT18), .A2(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n387), .A2(new_n391), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n330), .A2(G140), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n402), .A2(new_n414), .A3(KEYINPUT74), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT74), .B1(new_n402), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n195), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n398), .A2(new_n400), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n195), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n379), .B1(new_n409), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n395), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n422), .A2(new_n392), .A3(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n408), .A2(new_n407), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n379), .B(new_n420), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n280), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n429));
  INV_X1    g243(.A(new_n379), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n431), .B2(new_n425), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n434), .A3(G475), .ZN(new_n435));
  INV_X1    g249(.A(new_n406), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n415), .B2(new_n416), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n398), .A2(KEYINPUT19), .A3(new_n400), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n195), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n436), .B(new_n440), .C1(new_n422), .C2(new_n392), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n379), .B1(new_n441), .B2(new_n420), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n405), .B(new_n406), .C1(new_n392), .C2(KEYINPUT17), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n419), .A2(new_n413), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n443), .A2(new_n396), .B1(new_n444), .B2(new_n411), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n445), .B2(new_n379), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n280), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT20), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n441), .A2(new_n420), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n425), .B1(new_n450), .B2(new_n379), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n447), .A4(new_n280), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n435), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G116), .B(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(new_n206), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n197), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n230), .A2(G143), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT13), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G134), .C1(KEYINPUT13), .C2(new_n458), .ZN(new_n461));
  XNOR2_X1  g275(.A(G128), .B(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n239), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(KEYINPUT93), .A3(new_n239), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n457), .A2(new_n461), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n295), .A2(G122), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n206), .B1(new_n468), .B2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g283(.A(new_n456), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n458), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G134), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n463), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n456), .A2(new_n206), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G217), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n187), .A2(new_n477), .A3(G953), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n467), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n467), .B2(new_n476), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n280), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI221_X1 g298(.A(new_n280), .B1(KEYINPUT15), .B2(new_n482), .C1(new_n479), .C2(new_n480), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT94), .Z(new_n487));
  INV_X1    g301(.A(G952), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(G953), .ZN(new_n489));
  INV_X1    g303(.A(G234), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n280), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n455), .A2(new_n487), .A3(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n288), .A2(new_n376), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT26), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G101), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT68), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT68), .B1(new_n499), .B2(new_n501), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n382), .B2(G210), .ZN(new_n507));
  OAI211_X1 g321(.A(G210), .B(new_n191), .C1(new_n388), .C2(new_n389), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n382), .A2(new_n506), .A3(G210), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n504), .C2(new_n503), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n510), .B2(new_n513), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n519));
  XNOR2_X1  g333(.A(G134), .B(G137), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT64), .B1(new_n520), .B2(new_n246), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n241), .A2(G134), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n243), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT64), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(new_n247), .A3(new_n231), .A4(new_n229), .ZN(new_n527));
  INV_X1    g341(.A(new_n318), .ZN(new_n528));
  INV_X1    g342(.A(new_n203), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n248), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n519), .B(KEYINPUT28), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n524), .B1(new_n523), .B2(G131), .ZN(new_n538));
  AOI211_X1 g352(.A(KEYINPUT64), .B(new_n246), .C1(new_n522), .C2(new_n243), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n229), .A2(new_n247), .A3(new_n231), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n203), .B1(new_n247), .B2(new_n245), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n318), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n534), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n519), .B1(new_n545), .B2(KEYINPUT28), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n518), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT30), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n527), .A2(new_n549), .A3(new_n530), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n531), .B1(new_n551), .B2(new_n318), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n517), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT29), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n536), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(KEYINPUT28), .B2(new_n545), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT29), .A3(new_n518), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n280), .ZN(new_n558));
  OAI21_X1  g372(.A(G472), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n517), .B1(new_n537), .B2(new_n546), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT70), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n552), .B2(new_n518), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n528), .B1(new_n548), .B2(new_n550), .ZN(new_n564));
  NOR4_X1   g378(.A1(new_n564), .A2(new_n517), .A3(KEYINPUT31), .A4(new_n531), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(new_n517), .C1(new_n537), .C2(new_n546), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n559), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT76), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT71), .B1(new_n299), .B2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT23), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n299), .A2(G128), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n230), .A2(G119), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT71), .A3(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n578), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT24), .B(G110), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n584), .A2(KEYINPUT73), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT73), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n436), .B(new_n417), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n407), .ZN(new_n591));
  OAI221_X1 g405(.A(new_n591), .B1(new_n583), .B2(new_n582), .C1(new_n585), .C2(new_n586), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n597), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n477), .B1(G234), .B2(new_n280), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n280), .A3(new_n600), .ZN(new_n606));
  NOR2_X1   g420(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n574), .A2(new_n575), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n575), .B1(new_n574), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n498), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n569), .B2(new_n280), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n569), .A2(new_n614), .A3(new_n280), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n617), .A3(G472), .A4(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n569), .A2(new_n614), .A3(new_n280), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n620), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n569), .A2(new_n571), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n609), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n288), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n290), .B(new_n496), .C1(new_n358), .C2(new_n374), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n479), .A2(new_n480), .ZN(new_n632));
  AND2_X1   g446(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n632), .B1(new_n635), .B2(new_n633), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(G478), .A3(new_n280), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(KEYINPUT98), .A2(G478), .ZN(new_n638));
  AND2_X1   g452(.A1(KEYINPUT98), .A2(G478), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n481), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n435), .B2(new_n454), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AND2_X1   g462(.A1(new_n435), .A2(new_n454), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n630), .A2(new_n649), .A3(new_n487), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n629), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n206), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n608), .A2(new_n602), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT36), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n594), .B1(new_n656), .B2(new_n597), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n593), .A2(KEYINPUT36), .A3(new_n599), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n603), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n498), .A2(new_n625), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n574), .A2(new_n661), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n288), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT101), .B(G900), .Z(new_n667));
  AND2_X1   g481(.A1(new_n494), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n492), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n649), .A2(new_n487), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n376), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT103), .B(G128), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G30));
  INV_X1    g491(.A(new_n288), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n672), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n572), .A2(new_n573), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n552), .A2(new_n517), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n280), .B1(new_n518), .B2(new_n545), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n358), .A2(new_n374), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n455), .A2(new_n487), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n661), .A2(new_n290), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n681), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  INV_X1    g508(.A(new_n672), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n695), .B(new_n641), .C1(new_n435), .C2(new_n454), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n375), .A3(KEYINPUT104), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT104), .B1(new_n696), .B2(new_n375), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n666), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n284), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n275), .B1(new_n258), .B2(new_n262), .ZN(new_n705));
  OAI22_X1  g519(.A1(new_n273), .A2(new_n270), .B1(new_n705), .B2(new_n194), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n189), .B1(new_n706), .B2(new_n280), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n703), .B(new_n189), .C1(new_n706), .C2(new_n280), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n188), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n574), .A2(new_n609), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT106), .B(new_n188), .C1(new_n708), .C2(new_n709), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n714), .A3(new_n644), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n712), .A2(new_n714), .A3(new_n650), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  OAI211_X1 g534(.A(new_n188), .B(new_n375), .C1(new_n708), .C2(new_n709), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n721), .A2(new_n665), .A3(new_n497), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  OAI21_X1  g537(.A(new_n566), .B1(new_n518), .B2(new_n556), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n571), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n621), .B1(new_n569), .B2(new_n280), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g542(.A(KEYINPUT107), .B(new_n621), .C1(new_n569), .C2(new_n280), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n626), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n375), .A2(new_n689), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n496), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n712), .A2(new_n715), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT108), .B(G122), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G24));
  INV_X1    g549(.A(new_n721), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n728), .A2(new_n729), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT109), .B1(new_n737), .B2(new_n661), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n608), .A2(new_n602), .B1(new_n603), .B2(new_n659), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n728), .A2(new_n739), .A3(new_n729), .A4(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n696), .B(new_n736), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND3_X1  g557(.A1(new_n358), .A2(new_n289), .A3(new_n374), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n358), .A2(new_n374), .A3(KEYINPUT111), .A4(new_n289), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n746), .A2(new_n188), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n284), .A2(new_n286), .ZN(new_n750));
  INV_X1    g564(.A(new_n272), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n263), .A2(new_n277), .A3(new_n194), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n281), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n276), .A2(new_n277), .ZN(new_n754));
  OAI211_X1 g568(.A(G469), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n749), .A2(new_n755), .A3(new_n284), .A4(new_n286), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n758), .A3(KEYINPUT112), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n746), .A2(new_n188), .A3(new_n747), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n279), .B2(new_n287), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n749), .A3(new_n284), .A4(new_n286), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n713), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT42), .B1(new_n766), .B2(new_n696), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n696), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND2_X1  g585(.A1(new_n759), .A2(new_n765), .ZN(new_n772));
  INV_X1    g586(.A(new_n673), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n714), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  INV_X1    g589(.A(new_n284), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n274), .A2(new_n278), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n751), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n778), .A2(KEYINPUT113), .A3(KEYINPUT45), .A4(new_n751), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n189), .B1(new_n779), .B2(new_n780), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n286), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n776), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT46), .B(new_n286), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n711), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n679), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n746), .A2(new_n747), .ZN(new_n794));
  INV_X1    g608(.A(new_n625), .ZN(new_n795));
  INV_X1    g609(.A(new_n641), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n649), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT43), .Z(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n661), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n794), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  INV_X1    g618(.A(new_n696), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n794), .A2(new_n574), .A3(new_n805), .A4(new_n609), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n790), .A2(new_n791), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n807), .B2(new_n188), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n809), .B(new_n711), .C1(new_n790), .C2(new_n791), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n806), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n806), .C1(new_n808), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  NOR3_X1   g630(.A1(new_n761), .A2(new_n710), .A3(new_n492), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n798), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n714), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n798), .A2(new_n493), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n730), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n488), .B(G953), .C1(new_n823), .C2(new_n736), .ZN(new_n824));
  INV_X1    g638(.A(new_n686), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n817), .A2(new_n609), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n642), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n824), .A2(KEYINPUT122), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT122), .B1(new_n824), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n820), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n794), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n808), .A2(new_n810), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n710), .A2(new_n188), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OR4_X1    g650(.A1(new_n711), .A2(new_n688), .A3(new_n710), .A4(new_n289), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT121), .B1(new_n822), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n818), .B1(new_n738), .B2(new_n741), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n649), .A3(new_n641), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT51), .B1(new_n836), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n844), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n808), .A2(new_n810), .A3(new_n834), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n832), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n830), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n666), .B1(new_n699), .B2(new_n674), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n661), .A2(new_n711), .A3(new_n695), .ZN(new_n852));
  INV_X1    g666(.A(new_n731), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n758), .A2(new_n852), .A3(new_n686), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n742), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n742), .A2(new_n857), .A3(new_n851), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n484), .A2(KEYINPUT117), .A3(new_n485), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT117), .B1(new_n484), .B2(new_n485), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n863));
  OAI21_X1  g677(.A(G475), .B1(new_n432), .B2(new_n433), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n862), .B(new_n454), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n435), .A2(KEYINPUT118), .A3(new_n454), .A4(new_n862), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n496), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n375), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n375), .A2(new_n642), .A3(KEYINPUT116), .A4(new_n870), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT116), .B1(new_n630), .B2(new_n642), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n625), .B(new_n627), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n665), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n455), .A2(new_n695), .A3(new_n862), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n831), .A3(new_n678), .A4(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n612), .A2(new_n875), .A3(new_n662), .A4(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n726), .A2(new_n727), .ZN(new_n880));
  INV_X1    g694(.A(new_n729), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n725), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n740), .B1(new_n882), .B2(new_n739), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n661), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n805), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n772), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n879), .A2(new_n774), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n859), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n716), .A2(new_n719), .A3(new_n733), .A4(new_n722), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND4_X1   g704(.A1(KEYINPUT42), .A2(new_n772), .A3(new_n714), .A4(new_n696), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n767), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n893), .A3(KEYINPUT53), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n875), .A2(new_n878), .A3(new_n612), .A4(new_n662), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n885), .B2(new_n772), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n774), .A3(new_n856), .A4(new_n858), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(KEYINPUT119), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n774), .A4(new_n886), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n859), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n890), .C1(new_n891), .C2(new_n767), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n899), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n901), .A2(new_n902), .A3(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n908), .A2(new_n909), .A3(new_n899), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n894), .B2(new_n899), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT120), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n850), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n710), .B(KEYINPUT49), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n609), .A2(new_n188), .A3(new_n289), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n688), .A2(new_n797), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n919), .A3(new_n825), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(G75));
  XNOR2_X1  g735(.A(new_n366), .B(new_n347), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n280), .B1(new_n908), .B2(new_n899), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(G210), .ZN(new_n926));
  OR2_X1    g740(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n191), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n926), .A2(new_n924), .A3(new_n927), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n706), .B(KEYINPUT124), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n908), .A2(new_n899), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT54), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n910), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n285), .B(KEYINPUT57), .Z(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n786), .A2(new_n787), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n925), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n929), .B1(new_n940), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n925), .A2(new_n451), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n451), .B1(new_n925), .B2(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n929), .ZN(G60));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n634), .A2(new_n636), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n937), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n909), .B1(new_n908), .B2(new_n899), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n948), .B(new_n953), .C1(new_n912), .C2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n930), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n914), .A2(new_n911), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n950), .B1(new_n959), .B2(new_n952), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(G63));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n908), .A2(new_n899), .ZN(new_n963));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n601), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n908), .B2(new_n899), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n929), .B1(new_n967), .B2(new_n659), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n495), .B2(new_n333), .ZN(new_n972));
  AND4_X1   g786(.A1(new_n612), .A2(new_n890), .A3(new_n662), .A4(new_n875), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n355), .B(new_n356), .C1(G898), .C2(new_n191), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  NAND2_X1  g790(.A1(new_n438), .A2(new_n439), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n551), .B(new_n977), .Z(new_n978));
  NAND2_X1  g792(.A1(G900), .A2(G953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n802), .B1(new_n713), .B2(new_n731), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n792), .A3(new_n679), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n742), .A2(new_n851), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n774), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n770), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n814), .B2(new_n812), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n980), .B1(new_n986), .B2(new_n191), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n983), .A2(new_n693), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  INV_X1    g806(.A(new_n869), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n680), .B1(new_n993), .B2(new_n643), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n994), .B(new_n831), .C1(new_n611), .C2(new_n610), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n992), .A2(new_n803), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n996), .B2(new_n815), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n988), .B(new_n990), .C1(new_n997), .C2(new_n978), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n978), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n989), .B1(new_n999), .B2(new_n987), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(G72));
  XNOR2_X1  g815(.A(new_n553), .B(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n986), .A2(new_n973), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n683), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n996), .A2(new_n815), .A3(new_n973), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n1005), .ZN(new_n1009));
  AND4_X1   g823(.A1(new_n553), .A2(new_n900), .A3(new_n1007), .A4(new_n1005), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1006), .A2(new_n1009), .A3(new_n929), .A4(new_n1010), .ZN(G57));
endmodule


