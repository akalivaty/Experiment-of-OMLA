//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(G211gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n207), .B2(new_n208), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(new_n216), .B2(G141gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n218), .A3(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n228), .C1(new_n218), .C2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n221), .B1(new_n224), .B2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n225), .A2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n213), .A2(new_n214), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n211), .A2(new_n212), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n203), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n202), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n231), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n207), .A2(new_n208), .ZN(new_n245));
  INV_X1    g044(.A(new_n209), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n247), .B2(new_n210), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n242), .B(new_n244), .C1(new_n248), .C2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT81), .B(new_n203), .C1(new_n232), .C2(KEYINPUT3), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n238), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n202), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n241), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n241), .B2(new_n255), .ZN(new_n258));
  OAI21_X1  g057(.A(G78gat), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G22gat), .ZN(new_n261));
  INV_X1    g060(.A(G78gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n255), .A3(new_n256), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT31), .B(G50gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G106gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n259), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n259), .B2(new_n264), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G226gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT64), .B(G169gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT24), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n273), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n286), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(KEYINPUT24), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G169gat), .A3(G176gat), .ZN(new_n295));
  AND4_X1   g094(.A1(KEYINPUT25), .A2(new_n292), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n278), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n275), .A2(new_n276), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(KEYINPUT26), .B2(new_n277), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n302), .A2(new_n283), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT27), .B(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n298), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n272), .B1(new_n313), .B2(new_n203), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n289), .A2(new_n297), .B1(new_n303), .B2(new_n311), .ZN(new_n315));
  INV_X1    g114(.A(new_n272), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n238), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n315), .B2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n272), .ZN(new_n321));
  INV_X1    g120(.A(new_n238), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n330), .B1(new_n324), .B2(new_n326), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n336), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT74), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  INV_X1    g145(.A(G120gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT1), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(G113gat), .B2(G120gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G127gat), .B(G134gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n234), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n242), .A2(new_n244), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n353), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n234), .A2(new_n353), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n234), .A2(new_n353), .A3(KEYINPUT79), .A4(new_n361), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n236), .A2(new_n233), .ZN(new_n367));
  INV_X1    g166(.A(new_n353), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT4), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n358), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n242), .A2(KEYINPUT3), .A3(new_n244), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n353), .B1(new_n234), .B2(new_n214), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT77), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n360), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n236), .A2(new_n361), .A3(new_n353), .A4(new_n233), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n382), .A3(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n375), .B1(new_n371), .B2(new_n372), .ZN(new_n386));
  INV_X1    g185(.A(new_n376), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n344), .B1(new_n378), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n232), .B(new_n235), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n361), .B1(new_n391), .B2(new_n353), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n364), .A2(new_n365), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n357), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n387), .A2(new_n386), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n343), .B(new_n388), .C1(new_n396), .C2(new_n360), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT6), .B(new_n344), .C1(new_n378), .C2(new_n389), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n269), .B1(new_n339), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n280), .A2(new_n281), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n291), .A2(new_n404), .A3(new_n279), .A4(new_n278), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n296), .A2(new_n278), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n405), .A2(new_n273), .B1(new_n406), .B2(new_n291), .ZN(new_n407));
  AND4_X1   g206(.A1(new_n283), .A2(new_n302), .A3(new_n310), .A4(new_n308), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n353), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n298), .A2(new_n368), .A3(new_n312), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n271), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n403), .ZN(new_n416));
  AOI211_X1 g215(.A(new_n413), .B(new_n416), .C1(new_n409), .C2(new_n410), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT71), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n409), .A2(new_n413), .A3(new_n410), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(KEYINPUT32), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT69), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n422), .A2(new_n424), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n407), .A2(new_n408), .A3(new_n353), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n368), .B1(new_n298), .B2(new_n312), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n414), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n416), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n414), .A3(new_n403), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT69), .B1(new_n425), .B2(new_n426), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n419), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n426), .A2(new_n428), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n415), .A2(new_n417), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n435), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n418), .A4(new_n427), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n439), .A2(new_n444), .A3(KEYINPUT36), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT36), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n402), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n377), .A2(new_n384), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n358), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n357), .B(new_n354), .C1(new_n355), .C2(new_n353), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT39), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n357), .B1(new_n377), .B2(new_n384), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n451), .B(new_n343), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(KEYINPUT84), .A3(new_n458), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT84), .B1(new_n457), .B2(new_n458), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n390), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n329), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n336), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n463), .A2(new_n464), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n399), .A2(new_n400), .A3(new_n333), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n332), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n332), .A2(KEYINPUT85), .A3(new_n476), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n329), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n318), .A2(new_n323), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT38), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n324), .A2(KEYINPUT37), .A3(new_n326), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT85), .B1(new_n332), .B2(new_n476), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n478), .B(KEYINPUT37), .C1(new_n324), .C2(new_n326), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n330), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT38), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n269), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n448), .B1(new_n474), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n267), .A2(new_n268), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n439), .A2(new_n444), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n464), .B2(new_n473), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n401), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n399), .A2(new_n400), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n471), .A2(new_n492), .A3(new_n498), .A4(new_n493), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(new_n497), .B1(KEYINPUT35), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT87), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n446), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n439), .A2(new_n444), .A3(KEYINPUT36), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n492), .B1(new_n471), .B2(new_n498), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n469), .A2(new_n470), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n472), .B1(new_n508), .B2(new_n335), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n507), .A2(new_n509), .A3(new_n462), .ZN(new_n510));
  INV_X1    g309(.A(new_n489), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n330), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n401), .A2(new_n333), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n492), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n506), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n516));
  INV_X1    g315(.A(new_n494), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n497), .C1(new_n507), .C2(new_n509), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n524), .A2(G1gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n527), .A2(new_n528), .A3(G8gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(G43gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G50gat), .ZN(new_n536));
  INV_X1    g335(.A(G50gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(G43gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(G43gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(G50gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT90), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n549), .ZN(new_n552));
  OR3_X1    g351(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n556), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .A4(new_n539), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(KEYINPUT89), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n543), .ZN(new_n564));
  INV_X1    g363(.A(new_n542), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n533), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n531), .A2(new_n532), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n551), .A2(new_n558), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(KEYINPUT17), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n559), .A2(KEYINPUT17), .A3(new_n566), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n523), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT18), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT11), .B(G169gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT12), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n574), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n523), .B(KEYINPUT13), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n569), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n568), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n576), .A2(new_n581), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n575), .B2(KEYINPUT18), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n581), .B1(new_n591), .B2(new_n583), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n583), .A3(new_n588), .ZN(new_n595));
  INV_X1    g394(.A(new_n581), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT92), .B1(new_n597), .B2(new_n589), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n570), .A2(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n570), .A2(KEYINPUT17), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n602), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n567), .A2(new_n614), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n619), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT9), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G71gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n262), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n625), .ZN(new_n632));
  AND2_X1   g431(.A1(G57gat), .A2(G64gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(G57gat), .A2(G64gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n625), .A2(KEYINPUT95), .A3(new_n626), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n629), .A2(new_n632), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n625), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n640));
  NAND3_X1  g439(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n639), .A2(new_n631), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(G57gat), .A2(G64gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(G57gat), .A2(G64gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(G71gat), .A2(G78gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n640), .B1(new_n649), .B2(new_n641), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n637), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(KEYINPUT96), .B(new_n637), .C1(new_n646), .C2(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n533), .B1(new_n655), .B2(KEYINPUT21), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT21), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(G231gat), .A2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(G127gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  INV_X1    g465(.A(new_n656), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n222), .ZN(new_n671));
  XNOR2_X1  g470(.A(G183gat), .B(G211gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n665), .A2(new_n668), .A3(new_n673), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n623), .A2(new_n624), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n653), .A2(new_n654), .A3(new_n612), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n646), .A2(new_n650), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n605), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n604), .A3(new_n609), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n604), .A2(new_n609), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n681), .A3(new_n605), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n680), .A2(new_n637), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n678), .A2(new_n679), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n655), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G230gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n271), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n678), .B2(new_n686), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G120gat), .B(G148gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(G176gat), .B(G204gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n698), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(KEYINPUT98), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n704), .B(new_n700), .C1(new_n701), .C2(new_n694), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n522), .A2(new_n600), .A3(new_n677), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n401), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g509(.A1(new_n507), .A2(new_n509), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT16), .B(G8gat), .Z(new_n712));
  AND3_X1   g511(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n530), .B1(new_n708), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT42), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(KEYINPUT42), .B2(new_n713), .ZN(G1325gat));
  INV_X1    g515(.A(G15gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n708), .A2(new_n717), .A3(new_n493), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n708), .A2(new_n504), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(G1326gat));
  NAND2_X1  g519(.A1(new_n708), .A2(new_n269), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT43), .B(G22gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  NAND2_X1  g522(.A1(new_n675), .A2(new_n676), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n706), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n624), .A2(new_n623), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT99), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n522), .A2(new_n600), .A3(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(G29gat), .A3(new_n498), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT45), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n597), .A2(new_n589), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n491), .A2(new_n500), .A3(KEYINPUT87), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n516), .B1(new_n515), .B2(new_n520), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n726), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT44), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n738), .B(new_n726), .C1(new_n491), .C2(new_n500), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT100), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n515), .A2(new_n520), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT100), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n738), .A4(new_n726), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n733), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n498), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n747), .ZN(G1328gat));
  INV_X1    g547(.A(new_n711), .ZN(new_n749));
  OAI21_X1  g548(.A(G36gat), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n729), .A2(G36gat), .A3(new_n749), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(new_n493), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n729), .A2(G43gat), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n745), .A2(new_n504), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(G43gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g557(.A(new_n537), .B1(new_n745), .B2(new_n269), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n537), .B(new_n269), .C1(new_n729), .C2(KEYINPUT102), .ZN(new_n760));
  INV_X1    g559(.A(new_n728), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n599), .B(new_n761), .C1(new_n501), .C2(new_n521), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT48), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT103), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n733), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n740), .A2(new_n743), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n738), .B1(new_n522), .B2(new_n726), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n269), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G50gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT103), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n269), .A2(new_n537), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n762), .B2(new_n763), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n763), .B2(new_n762), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n771), .A2(new_n772), .A3(new_n775), .A4(KEYINPUT48), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n766), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT101), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n770), .A2(new_n778), .A3(G50gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n770), .B2(G50gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n760), .A2(new_n764), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n777), .B1(new_n782), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g582(.A(new_n732), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n677), .A2(new_n784), .A3(new_n706), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n741), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n401), .B(KEYINPUT104), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n711), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT49), .B(G64gat), .Z(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(G1333gat));
  NAND3_X1  g592(.A1(new_n786), .A2(G71gat), .A3(new_n504), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT105), .ZN(new_n795));
  INV_X1    g594(.A(new_n786), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n630), .B1(new_n796), .B2(new_n754), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n786), .A2(new_n269), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n724), .A2(new_n732), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n706), .B(new_n803), .C1(new_n768), .C2(new_n769), .ZN(new_n804));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804), .B2(new_n498), .ZN(new_n805));
  INV_X1    g604(.A(new_n726), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n515), .B2(new_n520), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n803), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n707), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n607), .A3(new_n401), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n805), .A2(new_n813), .ZN(G1336gat));
  NOR2_X1   g613(.A1(new_n804), .A2(new_n749), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n608), .ZN(new_n816));
  INV_X1    g615(.A(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n711), .A2(new_n608), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n821), .B1(new_n817), .B2(new_n818), .C1(new_n815), .C2(new_n608), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n804), .B2(new_n447), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n811), .ZN(new_n825));
  INV_X1    g624(.A(G99gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n754), .A2(new_n707), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(G1338gat));
  XOR2_X1   g628(.A(KEYINPUT107), .B(G106gat), .Z(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n804), .B2(new_n492), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n492), .A2(G106gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n812), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(G1339gat));
  NAND3_X1  g636(.A1(new_n677), .A2(new_n784), .A3(new_n707), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n601), .A2(new_n569), .A3(new_n602), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n523), .B1(new_n839), .B2(new_n568), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n568), .A2(new_n586), .A3(new_n585), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n580), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n589), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n698), .B1(new_n701), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n693), .A2(KEYINPUT54), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n689), .A2(new_n692), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT55), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n699), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n726), .A2(new_n843), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n843), .A2(KEYINPUT110), .A3(new_n706), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n589), .A2(new_n705), .A3(new_n703), .A4(new_n842), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n855), .B(new_n858), .C1(new_n784), .C2(new_n852), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n854), .B1(new_n859), .B2(new_n806), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n838), .B1(new_n860), .B2(new_n724), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT111), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(new_n838), .C1(new_n860), .C2(new_n724), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n787), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n495), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n732), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n865), .A2(new_n269), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n711), .A2(new_n498), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n754), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n599), .A2(new_n346), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1340gat));
  NOR4_X1   g675(.A1(new_n873), .A2(new_n347), .A3(new_n754), .A4(new_n707), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(new_n706), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n347), .ZN(G1341gat));
  INV_X1    g678(.A(new_n724), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n868), .A2(KEYINPUT112), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(G127gat), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT112), .B1(new_n868), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n880), .A2(new_n661), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(new_n874), .B2(new_n884), .ZN(G1342gat));
  INV_X1    g684(.A(G134gat), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n886), .A2(new_n867), .A3(new_n495), .A4(new_n726), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT56), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT113), .B(new_n886), .C1(new_n874), .C2(new_n726), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n726), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(G134gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(G1343gat));
  INV_X1    g692(.A(new_n872), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n504), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n492), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n856), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n706), .A2(KEYINPUT114), .A3(new_n589), .A4(new_n842), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n853), .B1(new_n594), .B2(new_n598), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT115), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n593), .B1(new_n590), .B2(new_n592), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n597), .A2(KEYINPUT92), .A3(new_n589), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n852), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n900), .A2(new_n901), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n806), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n854), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n904), .A2(new_n910), .A3(KEYINPUT116), .A4(new_n806), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n724), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT117), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n838), .B1(new_n915), .B2(KEYINPUT117), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n898), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n897), .B1(new_n865), .B2(new_n492), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n896), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n218), .B1(new_n921), .B2(new_n732), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n711), .A2(new_n492), .A3(new_n504), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n866), .A2(new_n787), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n600), .A2(new_n218), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT58), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n898), .ZN(new_n928));
  INV_X1    g727(.A(new_n838), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n912), .ZN(new_n930));
  INV_X1    g729(.A(new_n854), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n914), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n880), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n928), .B1(new_n935), .B2(new_n916), .ZN(new_n936));
  INV_X1    g735(.A(new_n920), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n600), .B(new_n895), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n924), .B2(new_n925), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT118), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n944), .B(new_n941), .C1(new_n938), .C2(G141gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n927), .B1(new_n943), .B2(new_n945), .ZN(G1344gat));
  AOI21_X1  g745(.A(new_n707), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n599), .A2(new_n677), .A3(new_n707), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n911), .A2(new_n931), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n948), .B(new_n950), .C1(new_n951), .C2(new_n724), .ZN(new_n952));
  INV_X1    g751(.A(new_n950), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n724), .B1(new_n911), .B2(new_n931), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n955), .A3(new_n269), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(new_n897), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n865), .A2(new_n928), .ZN(new_n958));
  OAI221_X1 g757(.A(new_n947), .B1(KEYINPUT120), .B2(new_n896), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n960));
  INV_X1    g759(.A(new_n924), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n707), .A2(G148gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(KEYINPUT119), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n964));
  INV_X1    g763(.A(new_n962), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n924), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n959), .A2(new_n960), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n216), .B1(new_n921), .B2(new_n706), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(KEYINPUT59), .B2(new_n968), .ZN(G1345gat));
  NOR3_X1   g768(.A1(new_n924), .A2(G155gat), .A3(new_n880), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n921), .A2(new_n724), .ZN(new_n972));
  OAI211_X1 g771(.A(KEYINPUT123), .B(new_n971), .C1(new_n972), .C2(new_n222), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n222), .B1(new_n921), .B2(new_n724), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1346gat));
  AOI21_X1  g776(.A(G162gat), .B1(new_n961), .B2(new_n726), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n806), .A2(new_n223), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n921), .B2(new_n979), .ZN(G1347gat));
  OR2_X1    g779(.A1(new_n749), .A2(new_n787), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n981), .A2(new_n754), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n871), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G169gat), .B1(new_n983), .B2(new_n599), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n865), .A2(new_n401), .A3(new_n749), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n517), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n784), .A2(new_n280), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1348gat));
  OAI21_X1  g787(.A(new_n276), .B1(new_n986), .B2(new_n707), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n706), .A2(G176gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g791(.A(G183gat), .B1(new_n983), .B2(new_n880), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n724), .A2(new_n304), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n986), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n983), .B2(new_n806), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT61), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n726), .A2(new_n305), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n986), .B2(new_n999), .ZN(G1351gat));
  NOR2_X1   g799(.A1(new_n504), .A2(new_n492), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(G197gat), .B1(new_n1003), .B2(new_n732), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n958), .B1(new_n897), .B2(new_n956), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n981), .A2(new_n504), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n600), .A2(G197gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1004), .B1(new_n1008), .B2(new_n1009), .ZN(G1352gat));
  XOR2_X1   g809(.A(KEYINPUT125), .B(G204gat), .Z(new_n1011));
  NAND2_X1  g810(.A1(new_n706), .A2(new_n1011), .ZN(new_n1012));
  OR3_X1    g811(.A1(new_n1002), .A2(KEYINPUT62), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g812(.A(KEYINPUT62), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n1005), .A2(new_n707), .A3(new_n1007), .ZN(new_n1015));
  OAI211_X1 g814(.A(new_n1013), .B(new_n1014), .C1(new_n1015), .C2(new_n1011), .ZN(G1353gat));
  NOR3_X1   g815(.A1(new_n1002), .A2(new_n204), .A3(new_n880), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n724), .B(new_n1006), .C1(new_n957), .C2(new_n958), .ZN(new_n1018));
  AOI21_X1  g817(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT63), .ZN(new_n1022));
  NOR3_X1   g821(.A1(new_n1005), .A2(new_n880), .A3(new_n1007), .ZN(new_n1023));
  INV_X1    g822(.A(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1025), .A2(KEYINPUT126), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1021), .A2(new_n1027), .ZN(G1354gat));
  INV_X1    g827(.A(G218gat), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1029), .B1(new_n1002), .B2(new_n806), .ZN(new_n1030));
  XNOR2_X1  g829(.A(new_n1030), .B(KEYINPUT127), .ZN(new_n1031));
  NOR2_X1   g830(.A1(new_n806), .A2(new_n1029), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1031), .B1(new_n1008), .B2(new_n1032), .ZN(G1355gat));
endmodule


