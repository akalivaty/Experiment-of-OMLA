//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G127gat), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n209), .A2(new_n217), .A3(KEYINPUT68), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT68), .B1(new_n209), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT23), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT64), .B(G169gat), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n224), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT24), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT25), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(KEYINPUT23), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT66), .B1(new_n242), .B2(new_n222), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n231), .A2(new_n233), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT24), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT25), .B1(new_n223), .B2(KEYINPUT23), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n236), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n222), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n238), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n239), .A2(new_n253), .A3(new_n241), .ZN(new_n254));
  INV_X1    g053(.A(new_n222), .ZN(new_n255));
  INV_X1    g054(.A(new_n223), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT26), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n235), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT27), .B(G183gat), .Z(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(G190gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n260), .A2(G190gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n259), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n221), .B1(new_n252), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n242), .A2(new_n222), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n234), .A2(new_n246), .A3(new_n236), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n251), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n228), .A2(new_n237), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n267), .A2(new_n262), .ZN(new_n281));
  INV_X1    g080(.A(new_n259), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n283), .A3(new_n220), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n271), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n294), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n284), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n271), .B1(new_n269), .B2(new_n284), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT71), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(KEYINPUT71), .A3(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(new_n270), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT34), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n305), .B1(new_n303), .B2(KEYINPUT71), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n297), .A3(new_n293), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G197gat), .ZN(new_n322));
  INV_X1    g121(.A(G197gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G204gat), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT73), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT73), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT22), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n325), .A2(new_n326), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n323), .A2(G204gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n321), .A2(G197gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n347));
  OAI21_X1  g146(.A(G218gat), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n332), .A3(new_n334), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n320), .B1(new_n351), .B2(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT79), .B1(new_n353), .B2(G141gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  INV_X1    g154(.A(G141gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(G148gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n356), .A3(G148gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n354), .A2(new_n357), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n362));
  INV_X1    g161(.A(G155gat), .ZN(new_n363));
  INV_X1    g162(.A(G162gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n353), .A2(G141gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n356), .A2(G148gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G155gat), .B(G162gat), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n319), .B1(new_n352), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n339), .A2(new_n350), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n336), .A2(new_n338), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n345), .A2(new_n349), .A3(new_n337), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT77), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n375), .B1(new_n339), .B2(new_n350), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n378), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n366), .A2(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n320), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n374), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n381), .A2(new_n383), .A3(new_n390), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n377), .B2(new_n378), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n373), .B1(new_n394), .B2(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT87), .B1(new_n396), .B2(new_n319), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398));
  INV_X1    g197(.A(new_n319), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n398), .B(new_n399), .C1(new_n393), .C2(new_n395), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n392), .B(new_n403), .C1(new_n397), .C2(new_n400), .ZN(new_n404));
  XOR2_X1   g203(.A(G78gat), .B(G106gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(KEYINPUT88), .A3(new_n404), .A4(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT88), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n411), .A2(new_n407), .B1(new_n402), .B2(new_n404), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n318), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n252), .B2(new_n268), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n381), .A2(new_n383), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(new_n280), .B2(new_n283), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n415), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n280), .B2(new_n283), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n389), .B1(new_n252), .B2(new_n268), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n422), .B2(new_n385), .ZN(new_n423));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n280), .A2(new_n283), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n415), .B1(new_n429), .B2(new_n389), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n384), .B(new_n380), .C1(new_n430), .C2(new_n420), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n419), .A3(new_n426), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n427), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n209), .A2(new_n217), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n386), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n373), .A2(new_n437), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT5), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n214), .A2(new_n216), .B1(new_n204), .B2(new_n206), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n209), .A2(new_n217), .A3(KEYINPUT68), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n373), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT82), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n386), .B1(new_n218), .B2(new_n219), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(new_n450), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n437), .B1(new_n386), .B2(new_n320), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n367), .A2(new_n320), .A3(new_n372), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(new_n387), .A3(KEYINPUT81), .A4(new_n437), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n457), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n443), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n442), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n438), .A2(new_n386), .A3(KEYINPUT4), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n469), .B(new_n470), .C1(new_n449), .C2(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n473), .A3(KEYINPUT85), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n465), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G57gat), .B(G85gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT84), .ZN(new_n477));
  XOR2_X1   g276(.A(G1gat), .B(G29gat), .Z(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n436), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(new_n475), .B2(new_n481), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n456), .A2(new_n464), .ZN(new_n484));
  INV_X1    g283(.A(new_n443), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n474), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT85), .B1(new_n464), .B2(new_n473), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n481), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT86), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n483), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n435), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n202), .B1(new_n413), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n411), .A2(new_n407), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n402), .A2(new_n404), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(new_n408), .A3(new_n317), .A4(new_n309), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n489), .B2(new_n490), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n475), .A2(new_n481), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n433), .A2(new_n434), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n493), .B(new_n432), .C1(new_n501), .C2(new_n502), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n419), .C1(new_n422), .C2(new_n385), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n431), .A2(KEYINPUT91), .A3(new_n510), .A4(new_n419), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n426), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(new_n509), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n416), .B1(new_n418), .B2(new_n415), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(new_n383), .A3(new_n381), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n422), .A2(new_n385), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(KEYINPUT37), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n518), .A2(new_n524), .A3(new_n427), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n508), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n452), .A2(new_n450), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n527), .A2(new_n470), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n442), .B1(new_n528), .B2(new_n467), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT89), .B(KEYINPUT39), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n441), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT39), .B1(new_n532), .B2(new_n457), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n531), .B(new_n481), .C1(new_n529), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n489), .A2(new_n490), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n529), .A2(new_n533), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT40), .A3(new_n481), .A4(new_n531), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n498), .B(new_n408), .C1(new_n540), .C2(new_n504), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n409), .A2(new_n412), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n309), .A2(new_n317), .A3(KEYINPUT36), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT36), .B1(new_n309), .B2(new_n317), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n494), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n495), .A2(new_n507), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT13), .Z(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(G1gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT16), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n554), .B2(G1gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n556), .A3(G8gat), .ZN(new_n557));
  INV_X1    g356(.A(G8gat), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n551), .B(new_n555), .C1(new_n552), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G50gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G43gat), .ZN(new_n562));
  INV_X1    g361(.A(G43gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G50gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT15), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT95), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n564), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g368(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n565), .A2(KEYINPUT95), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n566), .A2(new_n569), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(KEYINPUT94), .B2(new_n572), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n576), .A2(new_n577), .B1(G29gat), .B2(G36gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n565), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n578), .A2(new_n565), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(new_n575), .A3(new_n557), .A4(new_n559), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n549), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(KEYINPUT17), .A3(new_n575), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n557), .A2(new_n559), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n548), .A3(new_n580), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n587), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT93), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT11), .B(G169gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(KEYINPUT93), .A3(new_n603), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n609), .A3(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n589), .A2(new_n590), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n579), .A2(new_n621), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n620), .A2(new_n623), .B1(KEYINPUT101), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n625), .A2(KEYINPUT101), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n627), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n626), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G57gat), .B(G64gat), .Z(new_n638));
  INV_X1    g437(.A(KEYINPUT9), .ZN(new_n639));
  INV_X1    g438(.A(G71gat), .ZN(new_n640));
  INV_X1    g439(.A(G78gat), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G71gat), .B(G78gat), .Z(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n560), .B1(KEYINPUT21), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT99), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G183gat), .B(G211gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n654), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n637), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n614), .A2(KEYINPUT103), .A3(new_n615), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n652), .A2(new_n665), .A3(new_n618), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n619), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT102), .B1(new_n647), .B2(new_n619), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n664), .B(new_n667), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n621), .A3(KEYINPUT10), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n676));
  INV_X1    g475(.A(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT104), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n675), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n684), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND4_X1   g488(.A1(new_n547), .A2(new_n607), .A3(new_n663), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n492), .A2(new_n493), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n435), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G8gat), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n690), .A2(new_n435), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT42), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n695), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n697), .B2(new_n699), .ZN(new_n705));
  INV_X1    g504(.A(new_n703), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT106), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(G1325gat));
  INV_X1    g507(.A(new_n318), .ZN(new_n709));
  AOI21_X1  g508(.A(G15gat), .B1(new_n690), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n544), .A2(new_n545), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G15gat), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT108), .Z(new_n719));
  AOI21_X1  g518(.A(new_n710), .B1(new_n719), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g519(.A1(new_n498), .A2(new_n408), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n690), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(new_n637), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n515), .A2(new_n524), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n483), .A2(new_n537), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n493), .A4(new_n432), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n543), .B1(new_n504), .B2(new_n540), .C1(new_n729), .C2(new_n517), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n691), .A2(new_n504), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT36), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n318), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n309), .A2(new_n317), .A3(KEYINPUT36), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n731), .A2(new_n721), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT35), .B1(new_n731), .B2(new_n499), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n413), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n725), .B(new_n726), .C1(new_n736), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n547), .B2(new_n637), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n689), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n605), .A2(new_n606), .ZN(new_n745));
  INV_X1    g544(.A(new_n662), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT110), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n691), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n730), .A2(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n726), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n747), .ZN(new_n753));
  INV_X1    g552(.A(G29gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(new_n692), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n753), .A2(new_n758), .A3(new_n754), .A4(new_n692), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n756), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n750), .B1(new_n760), .B2(new_n761), .ZN(G1328gat));
  AOI21_X1  g561(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n753), .A2(new_n435), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G36gat), .B1(new_n749), .B2(new_n504), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1329gat));
  OAI21_X1  g567(.A(new_n725), .B1(new_n751), .B2(new_n726), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n547), .A2(KEYINPUT44), .A3(new_n637), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n769), .A2(new_n711), .A3(new_n770), .A4(new_n748), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n563), .B1(new_n771), .B2(KEYINPUT112), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n743), .A2(new_n773), .A3(new_n711), .A4(new_n748), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n752), .A2(new_n563), .A3(new_n709), .A4(new_n747), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n769), .A2(new_n717), .A3(new_n770), .A4(new_n748), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G43gat), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT47), .B1(new_n781), .B2(new_n776), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(KEYINPUT113), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n777), .B1(new_n772), .B2(new_n774), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n782), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1330gat));
  NAND3_X1  g587(.A1(new_n743), .A2(new_n721), .A3(new_n748), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G50gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT48), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n753), .A2(new_n561), .A3(new_n721), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n790), .B(new_n793), .C1(new_n791), .C2(KEYINPUT48), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1331gat));
  NAND3_X1  g596(.A1(new_n744), .A2(new_n745), .A3(new_n663), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n751), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n692), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g600(.A1(new_n751), .A2(new_n504), .A3(new_n798), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  AND2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(G1333gat));
  NAND3_X1  g605(.A1(new_n799), .A2(G71gat), .A3(new_n717), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT115), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n799), .A2(new_n709), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n640), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT50), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1334gat));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n721), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g616(.A1(new_n607), .A2(new_n746), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n547), .A2(new_n637), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n547), .A2(KEYINPUT51), .A3(new_n637), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n752), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n818), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n689), .A2(new_n691), .A3(G85gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n607), .A2(new_n689), .A3(new_n746), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n769), .A2(new_n770), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n769), .A2(KEYINPUT116), .A3(new_n770), .A4(new_n828), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n831), .A2(new_n692), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n833), .B2(new_n611), .ZN(G1336gat));
  NOR3_X1   g633(.A1(new_n689), .A2(G92gat), .A3(new_n504), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n824), .A2(new_n825), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g636(.A(G92gat), .B1(new_n829), .B2(new_n504), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n840), .A3(new_n823), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n819), .A2(KEYINPUT118), .A3(new_n820), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n841), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n831), .A2(new_n435), .A3(new_n832), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(G92gat), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n845), .B2(new_n837), .ZN(G1337gat));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n717), .A3(new_n832), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G99gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n689), .A2(new_n318), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(G99gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n824), .A2(new_n825), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(G1338gat));
  INV_X1    g652(.A(G106gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n744), .A2(new_n854), .A3(new_n721), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n824), .A2(new_n825), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858));
  OAI21_X1  g657(.A(G106gat), .B1(new_n829), .B2(new_n543), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n841), .A2(new_n842), .A3(new_n856), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n721), .A3(new_n832), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(G106gat), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n860), .B1(new_n863), .B2(new_n858), .ZN(G1339gat));
  NAND3_X1  g663(.A1(new_n663), .A2(new_n745), .A3(new_n689), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n582), .A2(new_n586), .A3(new_n549), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n548), .B1(new_n592), .B2(new_n580), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n602), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n587), .A2(new_n595), .A3(new_n596), .A4(new_n603), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n687), .B2(new_n688), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n675), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n677), .B1(new_n671), .B2(new_n672), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n685), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT55), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(KEYINPUT55), .A3(new_n877), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n605), .A2(new_n606), .A3(new_n686), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n872), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n881), .A2(new_n632), .A3(new_n636), .A4(new_n686), .ZN(new_n884));
  INV_X1    g683(.A(new_n878), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n879), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n883), .A2(new_n726), .B1(new_n871), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n865), .B1(new_n889), .B2(new_n746), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n692), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n413), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n504), .ZN(new_n893));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n607), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n890), .A2(new_n543), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n691), .A2(new_n435), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n318), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n745), .A2(new_n212), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1340gat));
  NOR3_X1   g699(.A1(new_n897), .A2(new_n210), .A3(new_n850), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n893), .A2(new_n744), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n210), .ZN(G1341gat));
  INV_X1    g702(.A(new_n898), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n205), .A3(new_n662), .ZN(new_n905));
  AND4_X1   g704(.A1(new_n504), .A2(new_n891), .A3(new_n413), .A4(new_n746), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(G127gat), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1342gat));
  NOR2_X1   g709(.A1(new_n726), .A2(new_n435), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n203), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT56), .ZN(new_n913));
  OAI21_X1  g712(.A(G134gat), .B1(new_n904), .B2(new_n726), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(KEYINPUT56), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G1343gat));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n712), .A2(new_n896), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n890), .B2(new_n721), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n721), .A2(KEYINPUT57), .ZN(new_n923));
  INV_X1    g722(.A(new_n888), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n870), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n881), .A2(new_n686), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n607), .A2(new_n926), .A3(new_n885), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n637), .B1(new_n927), .B2(new_n872), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n662), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(new_n865), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n607), .B(new_n919), .C1(new_n922), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n917), .B1(new_n931), .B2(G141gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n543), .B1(new_n713), .B2(new_n715), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n890), .A2(new_n692), .A3(new_n933), .A4(new_n504), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n607), .A2(new_n356), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n931), .B2(G141gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n932), .A2(new_n937), .A3(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n939));
  AOI221_X4 g738(.A(new_n936), .B1(new_n917), .B2(new_n939), .C1(new_n931), .C2(G141gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(G1344gat));
  NAND2_X1  g740(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n870), .B1(new_n888), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n928), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n865), .B1(new_n945), .B2(new_n746), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT57), .B1(new_n946), .B2(new_n721), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n890), .A2(new_n721), .A3(new_n921), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n744), .ZN(new_n950));
  OAI211_X1 g749(.A(KEYINPUT59), .B(G148gat), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n922), .A2(new_n930), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n952), .A2(KEYINPUT59), .A3(new_n950), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT59), .ZN(new_n954));
  INV_X1    g753(.A(new_n934), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n744), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n951), .B(new_n953), .C1(new_n956), .C2(G148gat), .ZN(G1345gat));
  NOR3_X1   g756(.A1(new_n934), .A2(G155gat), .A3(new_n662), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n952), .A2(new_n662), .A3(new_n918), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n363), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT125), .B(new_n959), .C1(new_n960), .C2(new_n363), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1346gat));
  NOR3_X1   g764(.A1(new_n952), .A2(new_n726), .A3(new_n918), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n891), .A2(new_n933), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n911), .A2(new_n364), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n966), .A2(new_n364), .B1(new_n967), .B2(new_n968), .ZN(G1347gat));
  AND2_X1   g768(.A1(new_n890), .A2(new_n691), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n499), .A2(new_n504), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n225), .A3(new_n607), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n692), .A2(new_n504), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(new_n318), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n895), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G169gat), .B1(new_n979), .B2(new_n745), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n975), .A2(new_n980), .ZN(G1348gat));
  INV_X1    g780(.A(G176gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n974), .A2(new_n982), .A3(new_n744), .ZN(new_n983));
  OAI21_X1  g782(.A(G176gat), .B1(new_n979), .B2(new_n689), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1349gat));
  NOR2_X1   g784(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n986));
  OAI21_X1  g785(.A(G183gat), .B1(new_n979), .B2(new_n662), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n746), .A2(new_n264), .A3(new_n265), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n970), .A2(new_n971), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(G1350gat));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n232), .A3(new_n637), .ZN(new_n993));
  OAI21_X1  g792(.A(G190gat), .B1(new_n979), .B2(new_n726), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  AND3_X1   g796(.A1(new_n970), .A2(new_n435), .A3(new_n933), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n607), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n949), .A2(new_n717), .A3(new_n977), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n745), .A2(new_n323), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(G1352gat));
  OR2_X1    g801(.A1(new_n947), .A2(new_n948), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n717), .A2(new_n977), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1003), .A2(new_n744), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(G204gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n998), .A2(new_n321), .A3(new_n744), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(G1353gat));
  NAND4_X1  g809(.A1(new_n998), .A2(new_n328), .A3(new_n329), .A4(new_n746), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n746), .B(new_n1004), .C1(new_n947), .C2(new_n948), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1012), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G1354gat));
  NAND3_X1  g814(.A1(new_n1003), .A2(new_n637), .A3(new_n1004), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(G218gat), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n327), .A3(new_n637), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(G1355gat));
endmodule


