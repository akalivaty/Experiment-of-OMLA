//key=1010101010101010101010101010101010101010101010101010101010101010


module locked_locked_c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, 
        G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, 
        G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, 
        G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, 
        G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, 
        G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, 
        G409, G405, G402, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, 
        KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, 
        KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, 
        KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, 
        KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, 
        KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, 
        KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, 
        KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, 
        KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, 
        KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, 
        KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, 
        KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, 
        KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, 
        KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, 
        KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, 
        KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, 
        KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, 
        KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, 
        KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, 
        KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, 
        KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, 
        KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, 
        KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60,
         KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55,
         KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50,
         KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45,
         KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40,
         KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35,
         KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30,
         KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25,
         KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20,
         KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15,
         KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9,
         KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3,
         KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126,
         KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121,
         KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116,
         KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111,
         KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106,
         KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101,
         KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96,
         KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91,
         KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86,
         KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81,
         KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76,
         KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71,
         KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66,
         KEYINPUT65, KEYINPUT64;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
         G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063;

  AND2_X1 U1027 ( .A1(n1030), .A2(n1897), .ZN(n1029) );
  BUF_X1 U1028 ( .A(n1245), .Z(n1010) );
  XOR2_X1 U1029 ( .A(KEYINPUT89), .B(n1815), .Z(n1950) );
  XNOR2_X1 U1030 ( .A(n1358), .B(n1357), .ZN(n1476) );
  INV_X1 U1031 ( .A(n1807), .ZN(n1501) );
  NAND2_X1 U1032 ( .A1(n1349), .A2(n1348), .ZN(n1392) );
  AND2_X2 U1033 ( .A1(n1622), .A2(G330), .ZN(n1484) );
  AND2_X2 U1034 ( .A1(n1056), .A2(n1252), .ZN(n1055) );
  NAND2_X1 U1035 ( .A1(n1682), .A2(n1484), .ZN(n1506) );
  NOR2_X1 U1036 ( .A1(n2034), .A2(n1380), .ZN(n1382) );
  NOR2_X4 U1037 ( .A1(n1232), .A2(n1231), .ZN(n1368) );
  INV_X2 U1038 ( .A(n1114), .ZN(n1411) );
  XNOR2_X2 U1039 ( .A(n1093), .B(KEYINPUT2), .ZN(n1114) );
  XNOR2_X1 U1040 ( .A(G375), .B(G378), .ZN(n2063) );
  INV_X1 U1041 ( .A(G33), .ZN(n1740) );
  INV_X1 U1042 ( .A(KEYINPUT66), .ZN(n1011) );
  NAND2_X1 U1043 ( .A1(n1032), .A2(n1017), .ZN(n1031) );
  AND2_X1 U1044 ( .A1(n1511), .A2(n1681), .ZN(n1072) );
  XNOR2_X1 U1045 ( .A(n1404), .B(n1837), .ZN(n1897) );
  NOR2_X1 U1046 ( .A1(n1808), .A2(n1832), .ZN(n1819) );
  OR2_X1 U1047 ( .A1(n1213), .A2(n1829), .ZN(n2055) );
  NAND2_X1 U1048 ( .A1(n1087), .A2(n1086), .ZN(n1379) );
  OR2_X1 U1049 ( .A1(n2010), .A2(n1501), .ZN(n1087) );
  NAND2_X1 U1050 ( .A1(n1473), .A2(n1472), .ZN(n1682) );
  NAND2_X1 U1051 ( .A1(n1279), .A2(n1278), .ZN(n1052) );
  NOR2_X1 U1052 ( .A1(n1812), .A2(n1218), .ZN(n1810) );
  NOR2_X2 U1053 ( .A1(n1500), .A2(n1309), .ZN(n1503) );
  NOR2_X1 U1054 ( .A1(n1809), .A2(n1163), .ZN(n1218) );
  OR2_X1 U1055 ( .A1(n1359), .A2(n1494), .ZN(n1533) );
  NOR2_X1 U1056 ( .A1(n1470), .A2(n1274), .ZN(n1275) );
  AND2_X1 U1057 ( .A1(n1020), .A2(n1267), .ZN(n1268) );
  NAND2_X1 U1058 ( .A1(n1241), .A2(n1240), .ZN(n1474) );
  NOR2_X1 U1059 ( .A1(n1192), .A2(n1092), .ZN(n1194) );
  NOR2_X1 U1060 ( .A1(n1283), .A2(n1226), .ZN(n1227) );
  NOR2_X1 U1061 ( .A1(n1283), .A2(n1255), .ZN(n1256) );
  XNOR2_X1 U1062 ( .A(KEYINPUT4), .B(n1099), .ZN(n1317) );
  NOR2_X1 U1063 ( .A1(n1223), .A2(n1222), .ZN(n1287) );
  NAND2_X2 U1064 ( .A1(n1060), .A2(G13), .ZN(n1313) );
  NAND2_X1 U1065 ( .A1(G33), .A2(n1405), .ZN(n1097) );
  NAND2_X1 U1066 ( .A1(n2020), .A2(G20), .ZN(n1104) );
  INV_X1 U1067 ( .A(G1), .ZN(n2020) );
  NAND2_X1 U1068 ( .A1(G13), .A2(G1), .ZN(n1093) );
  XNOR2_X1 U1069 ( .A(n1097), .B(n1096), .ZN(n1098) );
  NAND2_X1 U1070 ( .A1(n1098), .A2(n1114), .ZN(n1234) );
  AND2_X1 U1071 ( .A1(n1313), .A2(n1317), .ZN(n1251) );
  INV_X1 U1072 ( .A(n1317), .ZN(n1297) );
  INV_X1 U1073 ( .A(n1897), .ZN(n1462) );
  XNOR2_X1 U1074 ( .A(n1265), .B(n1011), .ZN(n1020) );
  NOR2_X1 U1075 ( .A1(n1970), .A2(n1969), .ZN(n1971) );
  AND2_X2 U1076 ( .A1(n1411), .A2(n1040), .ZN(n1016) );
  NAND2_X1 U1077 ( .A1(n1411), .A2(n1740), .ZN(n1041) );
  INV_X1 U1078 ( .A(n1117), .ZN(n1079) );
  NAND2_X1 U1079 ( .A1(n1730), .A2(n1023), .ZN(n1069) );
  INV_X1 U1080 ( .A(KEYINPUT8), .ZN(n1326) );
  AND2_X1 U1081 ( .A1(G1698), .A2(n1740), .ZN(n1040) );
  XNOR2_X1 U1082 ( .A(n1250), .B(KEYINPUT17), .ZN(n1054) );
  INV_X1 U1083 ( .A(KEYINPUT81), .ZN(n1070) );
  NAND2_X1 U1084 ( .A1(n1012), .A2(n1048), .ZN(n1047) );
  NAND2_X1 U1085 ( .A1(n1501), .A2(n1050), .ZN(n1048) );
  NAND2_X1 U1086 ( .A1(n1234), .A2(G20), .ZN(n1099) );
  NAND2_X1 U1087 ( .A1(n1079), .A2(n1085), .ZN(n1292) );
  INV_X1 U1088 ( .A(n1104), .ZN(n1060) );
  NAND2_X1 U1089 ( .A1(n1079), .A2(n1024), .ZN(n1281) );
  NAND2_X1 U1090 ( .A1(n1198), .A2(n1197), .ZN(n1215) );
  XNOR2_X1 U1091 ( .A(n1195), .B(KEYINPUT7), .ZN(n1198) );
  AND2_X1 U1092 ( .A1(n1120), .A2(n1119), .ZN(n1127) );
  XNOR2_X1 U1093 ( .A(n1802), .B(KEYINPUT39), .ZN(n1808) );
  XOR2_X1 U1094 ( .A(KEYINPUT40), .B(n1950), .Z(n1817) );
  NOR2_X1 U1095 ( .A1(n1396), .A2(n1395), .ZN(n1404) );
  NAND2_X1 U1096 ( .A1(n1063), .A2(n1015), .ZN(n1736) );
  AND2_X1 U1097 ( .A1(n1069), .A2(n1064), .ZN(n1063) );
  NAND2_X1 U1098 ( .A1(n1067), .A2(n1065), .ZN(n1064) );
  NAND2_X1 U1099 ( .A1(n1392), .A2(n1807), .ZN(n1028) );
  XNOR2_X1 U1100 ( .A(G384), .B(G396), .ZN(n1963) );
  XNOR2_X1 U1101 ( .A(n1486), .B(KEYINPUT52), .ZN(n1798) );
  NOR2_X1 U1102 ( .A1(n1027), .A2(G41), .ZN(n1026) );
  INV_X1 U1103 ( .A(G294), .ZN(n1027) );
  NAND2_X1 U1104 ( .A1(n1079), .A2(n1078), .ZN(n1247) );
  AND2_X1 U1105 ( .A1(G116), .A2(n1085), .ZN(n1078) );
  BUF_X1 U1106 ( .A(n1223), .Z(n1330) );
  NAND2_X1 U1107 ( .A1(n1411), .A2(G33), .ZN(n1117) );
  OR2_X1 U1108 ( .A1(n1292), .A2(n1082), .ZN(n1312) );
  INV_X1 U1109 ( .A(G97), .ZN(n1082) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(G41), .ZN(n1024) );
  OR2_X1 U1111 ( .A1(n1292), .A2(n1081), .ZN(n1173) );
  INV_X1 U1112 ( .A(G77), .ZN(n1081) );
  NOR2_X2 U1113 ( .A1(n1115), .A2(n1330), .ZN(n1196) );
  INV_X1 U1114 ( .A(G68), .ZN(n1084) );
  INV_X1 U1115 ( .A(KEYINPUT34), .ZN(n1153) );
  NAND2_X1 U1116 ( .A1(n1018), .A2(n1035), .ZN(n1034) );
  AND2_X1 U1117 ( .A1(n1037), .A2(n1036), .ZN(n1266) );
  OR2_X1 U1118 ( .A1(n1292), .A2(n1083), .ZN(n1101) );
  NAND2_X1 U1119 ( .A1(n2014), .A2(n1070), .ZN(n1066) );
  NAND2_X1 U1120 ( .A1(n1068), .A2(n1070), .ZN(n1067) );
  NAND2_X1 U1121 ( .A1(n2016), .A2(KEYINPUT81), .ZN(n1062) );
  OR2_X1 U1122 ( .A1(n1051), .A2(n1043), .ZN(n1042) );
  OR2_X1 U1123 ( .A1(n1501), .A2(n1050), .ZN(n1043) );
  AND2_X1 U1124 ( .A1(n1049), .A2(n1045), .ZN(n1044) );
  NAND2_X1 U1125 ( .A1(n1047), .A2(n1046), .ZN(n1045) );
  OR2_X1 U1126 ( .A1(n1012), .A2(n1022), .ZN(n1046) );
  NAND2_X1 U1127 ( .A1(n1200), .A2(n1199), .ZN(n1385) );
  OR2_X1 U1128 ( .A1(n1215), .A2(n1423), .ZN(n1199) );
  NAND2_X1 U1129 ( .A1(n1061), .A2(n1313), .ZN(n1059) );
  OR2_X1 U1130 ( .A1(n1861), .A2(G1), .ZN(n1061) );
  OR2_X1 U1131 ( .A1(n1292), .A2(n1025), .ZN(n1237) );
  NOR2_X1 U1132 ( .A1(n1495), .A2(n1497), .ZN(n1359) );
  NOR2_X1 U1133 ( .A1(n1289), .A2(n1288), .ZN(n1305) );
  INV_X1 U1134 ( .A(KEYINPUT92), .ZN(n1121) );
  NAND2_X1 U1135 ( .A1(n1385), .A2(n1383), .ZN(n1394) );
  XOR2_X1 U1136 ( .A(KEYINPUT29), .B(n1403), .Z(n1837) );
  AND2_X1 U1137 ( .A1(n1014), .A2(G330), .ZN(n1086) );
  INV_X1 U1138 ( .A(n1028), .ZN(n1467) );
  INV_X1 U1139 ( .A(KEYINPUT11), .ZN(n1357) );
  XNOR2_X1 U1140 ( .A(n1817), .B(n1816), .ZN(n1818) );
  INV_X1 U1141 ( .A(KEYINPUT90), .ZN(n1816) );
  XNOR2_X1 U1142 ( .A(n1484), .B(n1019), .ZN(n1485) );
  INV_X1 U1143 ( .A(KEYINPUT55), .ZN(n1071) );
  NOR2_X1 U1144 ( .A1(n1058), .A2(n2053), .ZN(n2054) );
  OR2_X1 U1145 ( .A1(n1494), .A2(n1807), .ZN(n1012) );
  AND2_X1 U1146 ( .A1(n1502), .A2(n2011), .ZN(n1013) );
  OR2_X1 U1147 ( .A1(n1378), .A2(n1807), .ZN(n1014) );
  OR2_X1 U1148 ( .A1(n1730), .A2(n1062), .ZN(n1015) );
  NOR2_X1 U1149 ( .A1(n1234), .A2(n1059), .ZN(n1245) );
  NAND2_X1 U1150 ( .A1(n1073), .A2(n1477), .ZN(n1622) );
  INV_X1 U1151 ( .A(G20), .ZN(n1085) );
  AND2_X1 U1152 ( .A1(n1087), .A2(n1014), .ZN(n1838) );
  OR2_X1 U1153 ( .A1(n1558), .A2(n1557), .ZN(n1017) );
  AND2_X1 U1154 ( .A1(n1334), .A2(n1091), .ZN(n1018) );
  NOR2_X1 U1155 ( .A1(n1343), .A2(n1342), .ZN(n1495) );
  AND2_X1 U1156 ( .A1(n1379), .A2(n1028), .ZN(n1730) );
  AND2_X1 U1157 ( .A1(n1483), .A2(n1482), .ZN(n1019) );
  AND2_X1 U1158 ( .A1(n1012), .A2(n1050), .ZN(n1021) );
  INV_X1 U1159 ( .A(G283), .ZN(n1025) );
  INV_X1 U1160 ( .A(G58), .ZN(n1083) );
  INV_X1 U1161 ( .A(G116), .ZN(n1080) );
  XNOR2_X1 U1162 ( .A(KEYINPUT114), .B(KEYINPUT53), .ZN(n1022) );
  AND2_X1 U1163 ( .A1(n1959), .A2(n1070), .ZN(n1023) );
  NOR2_X1 U1164 ( .A1(G41), .A2(n2002), .ZN(n2016) );
  NOR2_X2 U1165 ( .A1(G179), .A2(n1422), .ZN(n1937) );
  NOR2_X2 U1166 ( .A1(n1423), .A2(n1414), .ZN(n1921) );
  NAND2_X1 U1167 ( .A1(n1730), .A2(n1959), .ZN(n1469) );
  NAND2_X1 U1168 ( .A1(n1959), .A2(n1066), .ZN(n1065) );
  INV_X1 U1169 ( .A(n1959), .ZN(n1068) );
  NOR2_X2 U1170 ( .A1(n1423), .A2(n1422), .ZN(n1933) );
  NOR2_X2 U1171 ( .A1(G179), .A2(n1421), .ZN(n1922) );
  NOR2_X2 U1172 ( .A1(n1117), .A2(G41), .ZN(n1322) );
  NAND2_X1 U1173 ( .A1(n1079), .A2(n1026), .ZN(n1254) );
  XNOR2_X1 U1174 ( .A(n1029), .B(n1960), .ZN(n1898) );
  INV_X1 U1175 ( .A(n1822), .ZN(n1030) );
  XNOR2_X2 U1176 ( .A(n1031), .B(n1071), .ZN(G387) );
  NAND2_X1 U1177 ( .A1(n1033), .A2(n1072), .ZN(n1032) );
  XNOR2_X1 U1178 ( .A(n1489), .B(n1488), .ZN(n1033) );
  NOR2_X1 U1179 ( .A1(n1340), .A2(n1423), .ZN(n1341) );
  XNOR2_X2 U1180 ( .A(n1034), .B(KEYINPUT74), .ZN(n1340) );
  XNOR2_X1 U1181 ( .A(n1074), .B(n1326), .ZN(n1035) );
  NOR2_X2 U1182 ( .A1(n1264), .A2(n1263), .ZN(n1366) );
  INV_X1 U1183 ( .A(n1264), .ZN(n1036) );
  NOR2_X1 U1184 ( .A1(n1263), .A2(G179), .ZN(n1037) );
  NOR2_X1 U1185 ( .A1(n1366), .A2(G169), .ZN(n1265) );
  INV_X1 U1186 ( .A(n1038), .ZN(n1039) );
  NAND2_X1 U1187 ( .A1(n1038), .A2(n1481), .ZN(n1279) );
  XNOR2_X2 U1188 ( .A(n1276), .B(KEYINPUT0), .ZN(n1038) );
  NAND2_X1 U1189 ( .A1(n1361), .A2(n1038), .ZN(n1362) );
  NAND2_X1 U1190 ( .A1(n1038), .A2(n1471), .ZN(n1473) );
  XNOR2_X1 U1191 ( .A(n1485), .B(n1039), .ZN(n1731) );
  NOR2_X2 U1192 ( .A1(n1041), .A2(G1698), .ZN(n1323) );
  NOR2_X1 U1193 ( .A1(n1041), .A2(G20), .ZN(n1310) );
  NAND2_X1 U1194 ( .A1(n1044), .A2(n1042), .ZN(n1499) );
  NAND2_X1 U1195 ( .A1(n1051), .A2(n1021), .ZN(n1049) );
  INV_X1 U1196 ( .A(n1022), .ZN(n1050) );
  XNOR2_X1 U1197 ( .A(n1493), .B(n1492), .ZN(n1051) );
  NOR2_X1 U1198 ( .A1(n1826), .A2(n1212), .ZN(n1213) );
  NAND2_X1 U1199 ( .A1(n1052), .A2(n1503), .ZN(n1490) );
  NAND2_X1 U1200 ( .A1(n1052), .A2(n1339), .ZN(n1349) );
  NAND2_X1 U1201 ( .A1(n1052), .A2(n1807), .ZN(n2011) );
  XNOR2_X2 U1202 ( .A(n1053), .B(n1253), .ZN(n1271) );
  NAND2_X1 U1203 ( .A1(n1055), .A2(n1054), .ZN(n1053) );
  NAND2_X1 U1204 ( .A1(n1057), .A2(n1717), .ZN(n1056) );
  INV_X1 U1205 ( .A(n1251), .ZN(n1057) );
  INV_X1 U1206 ( .A(n1392), .ZN(n1058) );
  INV_X1 U1207 ( .A(n1313), .ZN(n1203) );
  XNOR2_X2 U1208 ( .A(KEYINPUT67), .B(G33), .ZN(n1861) );
  INV_X1 U1209 ( .A(n1730), .ZN(n2019) );
  NAND2_X1 U1210 ( .A1(n1476), .A2(n1475), .ZN(n1073) );
  NAND2_X1 U1211 ( .A1(n1325), .A2(n1324), .ZN(n1074) );
  NAND2_X1 U1212 ( .A1(n1075), .A2(n2016), .ZN(n1466) );
  XNOR2_X1 U1213 ( .A(n1462), .B(n1076), .ZN(n1075) );
  XNOR2_X1 U1214 ( .A(n1822), .B(n1077), .ZN(n1076) );
  INV_X1 U1215 ( .A(KEYINPUT46), .ZN(n1077) );
  XNOR2_X2 U1216 ( .A(n1382), .B(n1381), .ZN(n1822) );
  OR2_X1 U1217 ( .A1(n1292), .A2(n1084), .ZN(n1137) );
  BUF_X1 U1218 ( .A(n1271), .Z(n1470) );
  AND2_X1 U1219 ( .A1(n1322), .A2(G77), .ZN(n1088) );
  NAND2_X1 U1220 ( .A1(n1824), .A2(n1823), .ZN(n1089) );
  AND2_X1 U1221 ( .A1(n1844), .A2(n1681), .ZN(n1090) );
  NOR2_X1 U1222 ( .A1(n1333), .A2(n1332), .ZN(n1091) );
  XOR2_X1 U1223 ( .A(KEYINPUT6), .B(n1191), .Z(n1092) );
  INV_X1 U1224 ( .A(n1331), .ZN(n1332) );
  INV_X1 U1225 ( .A(KEYINPUT65), .ZN(n1259) );
  INV_X1 U1226 ( .A(KEYINPUT3), .ZN(n1096) );
  XNOR2_X1 U1227 ( .A(n1533), .B(KEYINPUT113), .ZN(n1492) );
  NAND2_X1 U1228 ( .A1(n1152), .A2(n1193), .ZN(n1158) );
  INV_X1 U1229 ( .A(KEYINPUT69), .ZN(n1253) );
  INV_X1 U1230 ( .A(KEYINPUT110), .ZN(n1468) );
  NOR2_X1 U1231 ( .A1(n1160), .A2(n1420), .ZN(n1159) );
  XNOR2_X1 U1232 ( .A(n1469), .B(n1468), .ZN(n1487) );
  XNOR2_X1 U1233 ( .A(n1131), .B(KEYINPUT37), .ZN(n1826) );
  XNOR2_X1 U1234 ( .A(n1964), .B(n1963), .ZN(n1965) );
  BUF_X1 U1235 ( .A(n1411), .Z(n2007) );
  NAND2_X1 U1236 ( .A1(n1466), .A2(n1465), .ZN(G381) );
  INV_X1 U1237 ( .A(G13), .ZN(n2031) );
  INV_X1 U1238 ( .A(G50), .ZN(n2026) );
  NAND2_X1 U1239 ( .A1(n1203), .A2(n2026), .ZN(n1095) );
  NAND2_X1 U1240 ( .A1(n1310), .A2(G150), .ZN(n1094) );
  NAND2_X1 U1241 ( .A1(n1095), .A2(n1094), .ZN(n1103) );
  OR2_X1 U1242 ( .A1(G58), .A2(G68), .ZN(n2052) );
  AND2_X2 U1243 ( .A1(G20), .A2(G1), .ZN(n1405) );
  NAND2_X1 U1244 ( .A1(n2052), .A2(n1297), .ZN(n1100) );
  NAND2_X1 U1245 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
  NOR2_X1 U1246 ( .A1(n1103), .A2(n1102), .ZN(n1107) );
  INV_X1 U1247 ( .A(n1234), .ZN(n1105) );
  NAND2_X1 U1248 ( .A1(n1105), .A2(n1104), .ZN(n1132) );
  NAND2_X1 U1249 ( .A1(n1317), .A2(n1132), .ZN(n1206) );
  NAND2_X1 U1250 ( .A1(G50), .A2(n1206), .ZN(n1106) );
  NAND2_X1 U1251 ( .A1(n1107), .A2(n1106), .ZN(n1825) );
  NOR2_X1 U1252 ( .A1(G41), .A2(G45), .ZN(n1108) );
  NOR2_X1 U1253 ( .A1(G1), .A2(n1108), .ZN(n1115) );
  NAND2_X1 U1254 ( .A1(n1115), .A2(G274), .ZN(n1193) );
  NAND2_X1 U1255 ( .A1(n1016), .A2(G223), .ZN(n1109) );
  NAND2_X1 U1256 ( .A1(n1193), .A2(n1109), .ZN(n1112) );
  BUF_X2 U1257 ( .A(n1323), .Z(n1258) );
  NAND2_X1 U1258 ( .A1(n1258), .A2(G222), .ZN(n1110) );
  XOR2_X1 U1259 ( .A(KEYINPUT36), .B(n1110), .Z(n1111) );
  NOR2_X1 U1260 ( .A1(n1112), .A2(n1111), .ZN(n1120) );
  AND2_X1 U1261 ( .A1(G41), .A2(G33), .ZN(n1113) );
  NOR2_X1 U1262 ( .A1(n1114), .A2(n1113), .ZN(n1223) );
  NAND2_X1 U1263 ( .A1(n1196), .A2(G226), .ZN(n1116) );
  XNOR2_X1 U1264 ( .A(KEYINPUT91), .B(n1116), .ZN(n1118) );
  NOR2_X1 U1265 ( .A1(n1118), .A2(n1088), .ZN(n1119) );
  INV_X1 U1266 ( .A(G200), .ZN(n1420) );
  NOR2_X1 U1267 ( .A1(n1127), .A2(n1420), .ZN(n1122) );
  XNOR2_X1 U1268 ( .A(n1122), .B(n1121), .ZN(n1124) );
  NAND2_X1 U1269 ( .A1(n1127), .A2(G190), .ZN(n1123) );
  NAND2_X1 U1270 ( .A1(n1124), .A2(n1123), .ZN(n1125) );
  NOR2_X1 U1271 ( .A1(n1825), .A2(n1125), .ZN(n1130) );
  INV_X1 U1272 ( .A(G179), .ZN(n1233) );
  NAND2_X1 U1273 ( .A1(n1127), .A2(n1233), .ZN(n1126) );
  NAND2_X1 U1274 ( .A1(n1126), .A2(n1825), .ZN(n1129) );
  NOR2_X1 U1275 ( .A1(G169), .A2(n1127), .ZN(n1128) );
  NOR2_X1 U1276 ( .A1(n1129), .A2(n1128), .ZN(n1829) );
  NOR2_X1 U1277 ( .A1(n1130), .A2(n1829), .ZN(n1131) );
  INV_X1 U1278 ( .A(n1132), .ZN(n1177) );
  NAND2_X1 U1279 ( .A1(G58), .A2(n1177), .ZN(n1141) );
  NAND2_X1 U1280 ( .A1(n1310), .A2(G159), .ZN(n1134) );
  NAND2_X1 U1281 ( .A1(n1203), .A2(n1083), .ZN(n1133) );
  NAND2_X1 U1282 ( .A1(n1134), .A2(n1133), .ZN(n1139) );
  NAND2_X1 U1283 ( .A1(G58), .A2(G68), .ZN(n1135) );
  NAND2_X1 U1284 ( .A1(n2052), .A2(n1135), .ZN(n1628) );
  NAND2_X1 U1285 ( .A1(n1628), .A2(n1297), .ZN(n1136) );
  NAND2_X1 U1286 ( .A1(n1137), .A2(n1136), .ZN(n1138) );
  NOR2_X1 U1287 ( .A1(n1139), .A2(n1138), .ZN(n1140) );
  NAND2_X1 U1288 ( .A1(n1141), .A2(n1140), .ZN(n1142) );
  XNOR2_X1 U1289 ( .A(n1142), .B(KEYINPUT30), .ZN(n1809) );
  NAND2_X1 U1290 ( .A1(n1016), .A2(G226), .ZN(n1143) );
  XNOR2_X1 U1291 ( .A(n1143), .B(KEYINPUT32), .ZN(n1145) );
  NAND2_X1 U1292 ( .A1(G223), .A2(n1258), .ZN(n1144) );
  NAND2_X1 U1293 ( .A1(n1145), .A2(n1144), .ZN(n1146) );
  XNOR2_X1 U1294 ( .A(n1146), .B(KEYINPUT33), .ZN(n1148) );
  NAND2_X1 U1295 ( .A1(G232), .A2(n1196), .ZN(n1147) );
  NAND2_X1 U1296 ( .A1(n1148), .A2(n1147), .ZN(n1151) );
  NAND2_X1 U1297 ( .A1(n1322), .A2(G87), .ZN(n1149) );
  XNOR2_X1 U1298 ( .A(KEYINPUT31), .B(n1149), .ZN(n1150) );
  NOR2_X1 U1299 ( .A1(n1151), .A2(n1150), .ZN(n1152) );
  XOR2_X1 U1300 ( .A(KEYINPUT75), .B(n1233), .Z(n1423) );
  NOR2_X1 U1301 ( .A1(n1158), .A2(n1423), .ZN(n1154) );
  XNOR2_X1 U1302 ( .A(n1154), .B(n1153), .ZN(n1156) );
  NAND2_X1 U1303 ( .A1(n1158), .A2(G169), .ZN(n1155) );
  NAND2_X1 U1304 ( .A1(n1156), .A2(n1155), .ZN(n1157) );
  NAND2_X1 U1305 ( .A1(n1809), .A2(n1157), .ZN(n1833) );
  INV_X1 U1306 ( .A(n1833), .ZN(n1812) );
  INV_X1 U1307 ( .A(n1158), .ZN(n1160) );
  XNOR2_X1 U1308 ( .A(n1159), .B(KEYINPUT35), .ZN(n1162) );
  NAND2_X1 U1309 ( .A1(n1160), .A2(G190), .ZN(n1161) );
  NAND2_X1 U1310 ( .A1(n1162), .A2(n1161), .ZN(n1163) );
  NAND2_X1 U1311 ( .A1(n1258), .A2(G226), .ZN(n1164) );
  NAND2_X1 U1312 ( .A1(n1193), .A2(n1164), .ZN(n1168) );
  NAND2_X1 U1313 ( .A1(n1196), .A2(G238), .ZN(n1166) );
  NAND2_X1 U1314 ( .A1(G232), .A2(n1016), .ZN(n1165) );
  NAND2_X1 U1315 ( .A1(n1166), .A2(n1165), .ZN(n1167) );
  NOR2_X1 U1316 ( .A1(n1168), .A2(n1167), .ZN(n1170) );
  NAND2_X1 U1317 ( .A1(n1322), .A2(G97), .ZN(n1169) );
  NAND2_X1 U1318 ( .A1(n1170), .A2(n1169), .ZN(n1183) );
  NOR2_X1 U1319 ( .A1(G179), .A2(n1183), .ZN(n1172) );
  INV_X1 U1320 ( .A(n1183), .ZN(n1181) );
  NOR2_X1 U1321 ( .A1(G169), .A2(n1181), .ZN(n1171) );
  NOR2_X1 U1322 ( .A1(n1172), .A2(n1171), .ZN(n1180) );
  NAND2_X1 U1323 ( .A1(G50), .A2(n1310), .ZN(n1174) );
  NAND2_X1 U1324 ( .A1(n1174), .A2(n1173), .ZN(n1176) );
  NOR2_X1 U1325 ( .A1(G68), .A2(n1251), .ZN(n1175) );
  NOR2_X1 U1326 ( .A1(n1176), .A2(n1175), .ZN(n1179) );
  NAND2_X1 U1327 ( .A1(n1177), .A2(G68), .ZN(n1178) );
  NAND2_X1 U1328 ( .A1(n1179), .A2(n1178), .ZN(n1397) );
  NAND2_X1 U1329 ( .A1(n1180), .A2(n1397), .ZN(n1805) );
  INV_X1 U1330 ( .A(n1805), .ZN(n1400) );
  NAND2_X1 U1331 ( .A1(G190), .A2(n1181), .ZN(n1182) );
  XNOR2_X1 U1332 ( .A(n1182), .B(KEYINPUT28), .ZN(n1186) );
  NAND2_X1 U1333 ( .A1(G200), .A2(n1183), .ZN(n1184) );
  XOR2_X1 U1334 ( .A(KEYINPUT27), .B(n1184), .Z(n1185) );
  NAND2_X1 U1335 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
  NOR2_X1 U1336 ( .A1(n1397), .A2(n1187), .ZN(n1188) );
  NOR2_X1 U1337 ( .A1(n1400), .A2(n1188), .ZN(n1398) );
  INV_X1 U1338 ( .A(n1398), .ZN(n1219) );
  NAND2_X1 U1339 ( .A1(n1322), .A2(G107), .ZN(n1190) );
  NAND2_X1 U1340 ( .A1(G232), .A2(n1258), .ZN(n1189) );
  NAND2_X1 U1341 ( .A1(n1190), .A2(n1189), .ZN(n1192) );
  NAND2_X1 U1342 ( .A1(G238), .A2(n1016), .ZN(n1191) );
  NAND2_X1 U1343 ( .A1(n1194), .A2(n1193), .ZN(n1195) );
  NAND2_X1 U1344 ( .A1(n1196), .A2(G244), .ZN(n1197) );
  NAND2_X1 U1345 ( .A1(G169), .A2(n1215), .ZN(n1200) );
  NAND2_X1 U1346 ( .A1(G58), .A2(n1310), .ZN(n1202) );
  INV_X1 U1347 ( .A(G87), .ZN(n1778) );
  XOR2_X1 U1348 ( .A(KEYINPUT77), .B(n1778), .Z(n1605) );
  OR2_X1 U1349 ( .A1(n1605), .A2(n1292), .ZN(n1201) );
  NAND2_X1 U1350 ( .A1(n1202), .A2(n1201), .ZN(n1205) );
  NOR2_X1 U1351 ( .A1(G77), .A2(n1313), .ZN(n1204) );
  NOR2_X1 U1352 ( .A1(n1205), .A2(n1204), .ZN(n1208) );
  NAND2_X1 U1353 ( .A1(G77), .A2(n1206), .ZN(n1207) );
  NAND2_X1 U1354 ( .A1(n1208), .A2(n1207), .ZN(n1383) );
  NOR2_X1 U1355 ( .A1(n1219), .A2(n1394), .ZN(n1209) );
  NOR2_X1 U1356 ( .A1(n1400), .A2(n1209), .ZN(n1210) );
  NOR2_X1 U1357 ( .A1(n1218), .A2(n1210), .ZN(n1211) );
  NOR2_X1 U1358 ( .A1(n1812), .A2(n1211), .ZN(n1212) );
  XNOR2_X1 U1359 ( .A(n2055), .B(KEYINPUT93), .ZN(n1352) );
  INV_X1 U1360 ( .A(G190), .ZN(n1409) );
  NOR2_X1 U1361 ( .A1(n1215), .A2(n1409), .ZN(n1214) );
  NOR2_X1 U1362 ( .A1(n1383), .A2(n1214), .ZN(n1217) );
  NAND2_X1 U1363 ( .A1(G200), .A2(n1215), .ZN(n1216) );
  NAND2_X1 U1364 ( .A1(n1217), .A2(n1216), .ZN(n1391) );
  NAND2_X1 U1365 ( .A1(n1394), .A2(n1391), .ZN(n1387) );
  NOR2_X1 U1366 ( .A1(n1219), .A2(n1826), .ZN(n1220) );
  NAND2_X1 U1367 ( .A1(n1810), .A2(n1220), .ZN(n1221) );
  NOR2_X2 U1368 ( .A1(n1387), .A2(n1221), .ZN(n2035) );
  NAND2_X1 U1369 ( .A1(G45), .A2(n2020), .ZN(n1327) );
  NOR2_X1 U1370 ( .A1(n1327), .A2(G41), .ZN(n1222) );
  NAND2_X1 U1371 ( .A1(G270), .A2(n1287), .ZN(n1224) );
  XNOR2_X1 U1372 ( .A(n1224), .B(KEYINPUT10), .ZN(n1228) );
  INV_X1 U1373 ( .A(n1327), .ZN(n1225) );
  NAND2_X1 U1374 ( .A1(G274), .A2(n1225), .ZN(n1331) );
  NOR2_X1 U1375 ( .A1(G41), .A2(n1331), .ZN(n1283) );
  AND2_X1 U1376 ( .A1(G257), .A2(n1258), .ZN(n1226) );
  NAND2_X1 U1377 ( .A1(n1228), .A2(n1227), .ZN(n1232) );
  NAND2_X1 U1378 ( .A1(n1322), .A2(G303), .ZN(n1230) );
  NAND2_X1 U1379 ( .A1(n1016), .A2(G264), .ZN(n1229) );
  NAND2_X1 U1380 ( .A1(n1230), .A2(n1229), .ZN(n1231) );
  NAND2_X1 U1381 ( .A1(n1368), .A2(n1233), .ZN(n1242) );
  OR2_X1 U1382 ( .A1(n1010), .A2(n1297), .ZN(n1235) );
  NAND2_X1 U1383 ( .A1(n1235), .A2(G116), .ZN(n1241) );
  NAND2_X1 U1384 ( .A1(G97), .A2(n1310), .ZN(n1236) );
  NAND2_X1 U1385 ( .A1(n1237), .A2(n1236), .ZN(n1239) );
  NOR2_X1 U1386 ( .A1(G116), .A2(n1313), .ZN(n1238) );
  NOR2_X1 U1387 ( .A1(n1239), .A2(n1238), .ZN(n1240) );
  NAND2_X1 U1388 ( .A1(n1242), .A2(n1474), .ZN(n1244) );
  NOR2_X1 U1389 ( .A1(G169), .A2(n1368), .ZN(n1243) );
  NOR2_X1 U1390 ( .A1(n1244), .A2(n1243), .ZN(n1481) );
  NAND2_X1 U1391 ( .A1(G87), .A2(n1310), .ZN(n1252) );
  NAND2_X1 U1392 ( .A1(n1010), .A2(G107), .ZN(n1246) );
  XNOR2_X1 U1393 ( .A(n1246), .B(KEYINPUT68), .ZN(n1249) );
  XNOR2_X1 U1394 ( .A(KEYINPUT16), .B(n1247), .ZN(n1248) );
  NAND2_X1 U1395 ( .A1(n1249), .A2(n1248), .ZN(n1250) );
  XNOR2_X1 U1396 ( .A(n1254), .B(KEYINPUT14), .ZN(n1257) );
  AND2_X1 U1397 ( .A1(G257), .A2(n1016), .ZN(n1255) );
  NAND2_X1 U1398 ( .A1(n1257), .A2(n1256), .ZN(n1264) );
  NAND2_X1 U1399 ( .A1(n1258), .A2(G250), .ZN(n1262) );
  NAND2_X1 U1400 ( .A1(n1287), .A2(G264), .ZN(n1260) );
  XNOR2_X1 U1401 ( .A(n1260), .B(n1259), .ZN(n1261) );
  NAND2_X1 U1402 ( .A1(n1262), .A2(n1261), .ZN(n1263) );
  XNOR2_X1 U1403 ( .A(n1266), .B(KEYINPUT15), .ZN(n1267) );
  NAND2_X1 U1404 ( .A1(n1271), .A2(n1268), .ZN(n1270) );
  INV_X1 U1405 ( .A(KEYINPUT70), .ZN(n1269) );
  XNOR2_X2 U1406 ( .A(n1270), .B(n1269), .ZN(n1277) );
  INV_X1 U1407 ( .A(n1366), .ZN(n1372) );
  NAND2_X1 U1408 ( .A1(G200), .A2(n1372), .ZN(n1273) );
  NAND2_X1 U1409 ( .A1(G190), .A2(n1366), .ZN(n1272) );
  NAND2_X1 U1410 ( .A1(n1273), .A2(n1272), .ZN(n1274) );
  NOR2_X2 U1411 ( .A1(n1277), .A2(n1275), .ZN(n1276) );
  INV_X1 U1412 ( .A(n1277), .ZN(n1278) );
  NAND2_X1 U1413 ( .A1(n1323), .A2(G244), .ZN(n1280) );
  NAND2_X1 U1414 ( .A1(n1281), .A2(n1280), .ZN(n1282) );
  NOR2_X1 U1415 ( .A1(n1283), .A2(n1282), .ZN(n1285) );
  NAND2_X1 U1416 ( .A1(n1016), .A2(G250), .ZN(n1284) );
  NAND2_X1 U1417 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
  XNOR2_X1 U1418 ( .A(n1286), .B(KEYINPUT12), .ZN(n1289) );
  AND2_X1 U1419 ( .A1(G257), .A2(n1287), .ZN(n1288) );
  NOR2_X1 U1420 ( .A1(G169), .A2(n1305), .ZN(n1291) );
  INV_X1 U1421 ( .A(n1305), .ZN(n1369) );
  NOR2_X1 U1422 ( .A1(G179), .A2(n1369), .ZN(n1290) );
  NOR2_X1 U1423 ( .A1(n1291), .A2(n1290), .ZN(n1304) );
  NOR2_X1 U1424 ( .A1(G97), .A2(n1313), .ZN(n1294) );
  INV_X1 U1425 ( .A(G107), .ZN(n1717) );
  NOR2_X1 U1426 ( .A1(n1292), .A2(n1717), .ZN(n1293) );
  NOR2_X1 U1427 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
  XOR2_X1 U1428 ( .A(n1295), .B(KEYINPUT71), .Z(n1296) );
  XNOR2_X1 U1429 ( .A(KEYINPUT13), .B(n1296), .ZN(n1301) );
  NAND2_X1 U1430 ( .A1(n1310), .A2(G77), .ZN(n1299) );
  XOR2_X1 U1431 ( .A(n1717), .B(G97), .Z(n2023) );
  NAND2_X1 U1432 ( .A1(n2023), .A2(n1297), .ZN(n1298) );
  NAND2_X1 U1433 ( .A1(n1299), .A2(n1298), .ZN(n1300) );
  NOR2_X1 U1434 ( .A1(n1301), .A2(n1300), .ZN(n1303) );
  NAND2_X1 U1435 ( .A1(n1010), .A2(G97), .ZN(n1302) );
  NAND2_X1 U1436 ( .A1(n1303), .A2(n1302), .ZN(n1479) );
  NAND2_X1 U1437 ( .A1(n1304), .A2(n1479), .ZN(n1491) );
  INV_X1 U1438 ( .A(n1491), .ZN(n1500) );
  NAND2_X1 U1439 ( .A1(G200), .A2(n1369), .ZN(n1307) );
  NAND2_X1 U1440 ( .A1(G190), .A2(n1305), .ZN(n1306) );
  NAND2_X1 U1441 ( .A1(n1307), .A2(n1306), .ZN(n1308) );
  NOR2_X1 U1442 ( .A1(n1479), .A2(n1308), .ZN(n1309) );
  NAND2_X1 U1443 ( .A1(G68), .A2(n1310), .ZN(n1311) );
  NAND2_X1 U1444 ( .A1(n1312), .A2(n1311), .ZN(n1315) );
  NOR2_X1 U1445 ( .A1(G87), .A2(n1313), .ZN(n1314) );
  NOR2_X1 U1446 ( .A1(n1315), .A2(n1314), .ZN(n1321) );
  NAND2_X1 U1447 ( .A1(G87), .A2(n1010), .ZN(n1316) );
  NAND2_X1 U1448 ( .A1(n1317), .A2(n1316), .ZN(n1318) );
  NOR2_X1 U1449 ( .A1(G107), .A2(G97), .ZN(n1604) );
  NAND2_X1 U1450 ( .A1(n1604), .A2(n1605), .ZN(n1705) );
  NAND2_X1 U1451 ( .A1(n1318), .A2(n1705), .ZN(n1319) );
  XOR2_X1 U1452 ( .A(KEYINPUT9), .B(n1319), .Z(n1320) );
  NAND2_X1 U1453 ( .A1(n1321), .A2(n1320), .ZN(n1344) );
  NAND2_X1 U1454 ( .A1(n1322), .A2(G116), .ZN(n1334) );
  NAND2_X1 U1455 ( .A1(G244), .A2(n1016), .ZN(n1325) );
  NAND2_X1 U1456 ( .A1(n1323), .A2(G238), .ZN(n1324) );
  NAND2_X1 U1457 ( .A1(G250), .A2(n1327), .ZN(n1328) );
  XOR2_X1 U1458 ( .A(KEYINPUT73), .B(n1328), .Z(n1329) );
  NOR2_X1 U1459 ( .A1(n1330), .A2(n1329), .ZN(n1333) );
  INV_X1 U1460 ( .A(n1340), .ZN(n1363) );
  NAND2_X1 U1461 ( .A1(G190), .A2(n1363), .ZN(n1336) );
  NAND2_X1 U1462 ( .A1(G200), .A2(n1340), .ZN(n1335) );
  NAND2_X1 U1463 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
  NOR2_X1 U1464 ( .A1(n1344), .A2(n1337), .ZN(n1494) );
  XNOR2_X1 U1465 ( .A(n1494), .B(KEYINPUT78), .ZN(n1347) );
  INV_X1 U1466 ( .A(n1347), .ZN(n1338) );
  AND2_X1 U1467 ( .A1(n1503), .A2(n1338), .ZN(n1339) );
  XNOR2_X1 U1468 ( .A(n1341), .B(KEYINPUT76), .ZN(n1343) );
  INV_X1 U1469 ( .A(G169), .ZN(n1412) );
  NOR2_X1 U1470 ( .A1(n1412), .A2(n1363), .ZN(n1342) );
  INV_X1 U1471 ( .A(n1344), .ZN(n1497) );
  INV_X1 U1472 ( .A(n1359), .ZN(n1345) );
  AND2_X1 U1473 ( .A1(n1491), .A2(n1345), .ZN(n1346) );
  OR2_X1 U1474 ( .A1(n1347), .A2(n1346), .ZN(n1348) );
  NOR2_X1 U1475 ( .A1(G20), .A2(n2031), .ZN(n1406) );
  NAND2_X1 U1476 ( .A1(G213), .A2(n1406), .ZN(n1350) );
  NOR2_X1 U1477 ( .A1(G1), .A2(n1350), .ZN(n1834) );
  NAND2_X1 U1478 ( .A1(G343), .A2(n1834), .ZN(n1807) );
  NAND2_X1 U1479 ( .A1(n2035), .A2(n1467), .ZN(n1351) );
  NAND2_X1 U1480 ( .A1(n1352), .A2(n1351), .ZN(n2034) );
  INV_X1 U1481 ( .A(n1368), .ZN(n1375) );
  NAND2_X1 U1482 ( .A1(G200), .A2(n1375), .ZN(n1354) );
  NAND2_X1 U1483 ( .A1(G190), .A2(n1368), .ZN(n1353) );
  NAND2_X1 U1484 ( .A1(n1354), .A2(n1353), .ZN(n1355) );
  NOR2_X1 U1485 ( .A1(n1474), .A2(n1355), .ZN(n1356) );
  NOR2_X1 U1486 ( .A1(n1481), .A2(n1356), .ZN(n1358) );
  INV_X1 U1487 ( .A(n1476), .ZN(n1360) );
  NOR2_X1 U1488 ( .A1(n1360), .A2(n1533), .ZN(n1361) );
  INV_X1 U1489 ( .A(n1503), .ZN(n1478) );
  NOR2_X1 U1490 ( .A1(n1362), .A2(n1478), .ZN(n2010) );
  NOR2_X1 U1491 ( .A1(G179), .A2(n1363), .ZN(n1364) );
  NAND2_X1 U1492 ( .A1(n1369), .A2(n1364), .ZN(n1365) );
  NOR2_X1 U1493 ( .A1(n1366), .A2(n1365), .ZN(n1367) );
  NOR2_X1 U1494 ( .A1(n1368), .A2(n1367), .ZN(n1377) );
  NOR2_X1 U1495 ( .A1(n1340), .A2(n1369), .ZN(n1370) );
  XNOR2_X1 U1496 ( .A(KEYINPUT18), .B(n1370), .ZN(n1371) );
  NAND2_X1 U1497 ( .A1(n1371), .A2(G179), .ZN(n1373) );
  NOR2_X1 U1498 ( .A1(n1373), .A2(n1372), .ZN(n1374) );
  NOR2_X1 U1499 ( .A1(n1375), .A2(n1374), .ZN(n1376) );
  NOR2_X1 U1500 ( .A1(n1377), .A2(n1376), .ZN(n1378) );
  INV_X1 U1501 ( .A(n2035), .ZN(n2053) );
  NOR2_X1 U1502 ( .A1(n1379), .A2(n2053), .ZN(n1380) );
  INV_X1 U1503 ( .A(KEYINPUT38), .ZN(n1381) );
  NAND2_X1 U1504 ( .A1(n1383), .A2(n1501), .ZN(n1384) );
  XOR2_X1 U1505 ( .A(KEYINPUT5), .B(n1384), .Z(n1386) );
  NOR2_X1 U1506 ( .A1(n1385), .A2(n1386), .ZN(n1389) );
  AND2_X1 U1507 ( .A1(n1387), .A2(n1386), .ZN(n1388) );
  NOR2_X1 U1508 ( .A1(n1389), .A2(n1388), .ZN(n1839) );
  INV_X1 U1509 ( .A(n1839), .ZN(n1390) );
  NOR2_X2 U1510 ( .A1(n1379), .A2(n1390), .ZN(n1801) );
  XNOR2_X1 U1511 ( .A(n1801), .B(KEYINPUT88), .ZN(n1396) );
  NAND2_X1 U1512 ( .A1(n1392), .A2(n1391), .ZN(n1393) );
  NAND2_X1 U1513 ( .A1(n1394), .A2(n1393), .ZN(n1803) );
  AND2_X1 U1514 ( .A1(n1807), .A2(n1803), .ZN(n1395) );
  NAND2_X1 U1515 ( .A1(n1397), .A2(n1501), .ZN(n1399) );
  NAND2_X1 U1516 ( .A1(n1399), .A2(n1398), .ZN(n1402) );
  NAND2_X1 U1517 ( .A1(n1400), .A2(n1501), .ZN(n1401) );
  NAND2_X1 U1518 ( .A1(n1402), .A2(n1401), .ZN(n1403) );
  NAND2_X1 U1519 ( .A1(n1405), .A2(n2031), .ZN(n2002) );
  INV_X1 U1520 ( .A(n2016), .ZN(n2014) );
  NAND2_X1 U1521 ( .A1(n1406), .A2(G45), .ZN(n1407) );
  NAND2_X1 U1522 ( .A1(G1), .A2(n1407), .ZN(n1408) );
  XNOR2_X1 U1523 ( .A(KEYINPUT1), .B(n1408), .ZN(n1959) );
  NAND2_X1 U1524 ( .A1(n2014), .A2(n1959), .ZN(n1681) );
  NOR2_X1 U1525 ( .A1(n1085), .A2(G190), .ZN(n1427) );
  NAND2_X1 U1526 ( .A1(G200), .A2(n1427), .ZN(n1414) );
  NOR2_X1 U1527 ( .A1(G179), .A2(n1414), .ZN(n1934) );
  NAND2_X1 U1528 ( .A1(G77), .A2(n1934), .ZN(n1527) );
  NOR2_X1 U1529 ( .A1(n1085), .A2(n1409), .ZN(n1418) );
  NAND2_X1 U1530 ( .A1(G200), .A2(n1418), .ZN(n1422) );
  NAND2_X1 U1531 ( .A1(G97), .A2(n1937), .ZN(n1410) );
  NAND2_X1 U1532 ( .A1(n1527), .A2(n1410), .ZN(n1436) );
  NAND2_X1 U1533 ( .A1(G20), .A2(n1412), .ZN(n1413) );
  NAND2_X1 U1534 ( .A1(n2007), .A2(n1413), .ZN(n1884) );
  NOR2_X1 U1535 ( .A1(n1740), .A2(n1884), .ZN(n1909) );
  NAND2_X1 U1536 ( .A1(G116), .A2(n1921), .ZN(n1415) );
  NAND2_X1 U1537 ( .A1(n1909), .A2(n1415), .ZN(n1433) );
  AND2_X1 U1538 ( .A1(n1423), .A2(n1420), .ZN(n1416) );
  NAND2_X1 U1539 ( .A1(G190), .A2(n1416), .ZN(n1417) );
  NAND2_X1 U1540 ( .A1(G20), .A2(n1417), .ZN(n1928) );
  INV_X1 U1541 ( .A(n1928), .ZN(n1537) );
  NOR2_X1 U1542 ( .A1(n1537), .A2(n1778), .ZN(n1670) );
  NOR2_X1 U1543 ( .A1(n1423), .A2(G200), .ZN(n1426) );
  NAND2_X1 U1544 ( .A1(n1418), .A2(n1426), .ZN(n1654) );
  INV_X1 U1545 ( .A(n1654), .ZN(n1927) );
  AND2_X1 U1546 ( .A1(n1927), .A2(G283), .ZN(n1419) );
  NOR2_X1 U1547 ( .A1(n1670), .A2(n1419), .ZN(n1431) );
  NAND2_X1 U1548 ( .A1(n1427), .A2(n1420), .ZN(n1421) );
  NAND2_X1 U1549 ( .A1(n1922), .A2(G303), .ZN(n1425) );
  NAND2_X1 U1550 ( .A1(n1933), .A2(G294), .ZN(n1424) );
  NAND2_X1 U1551 ( .A1(n1425), .A2(n1424), .ZN(n1429) );
  NAND2_X1 U1552 ( .A1(n1427), .A2(n1426), .ZN(n1446) );
  NOR2_X1 U1553 ( .A1(n1717), .A2(n1446), .ZN(n1428) );
  NOR2_X1 U1554 ( .A1(n1429), .A2(n1428), .ZN(n1430) );
  NAND2_X1 U1555 ( .A1(n1431), .A2(n1430), .ZN(n1432) );
  NOR2_X1 U1556 ( .A1(n1433), .A2(n1432), .ZN(n1434) );
  XNOR2_X1 U1557 ( .A(n1434), .B(KEYINPUT103), .ZN(n1435) );
  NOR2_X1 U1558 ( .A1(n1436), .A2(n1435), .ZN(n1438) );
  NAND2_X1 U1559 ( .A1(n2031), .A2(n1861), .ZN(n1949) );
  NAND2_X1 U1560 ( .A1(n1949), .A2(n1884), .ZN(n1899) );
  NOR2_X1 U1561 ( .A1(G68), .A2(n1899), .ZN(n1437) );
  NOR2_X1 U1562 ( .A1(n1438), .A2(n1437), .ZN(n1457) );
  NAND2_X1 U1563 ( .A1(G128), .A2(n1922), .ZN(n1440) );
  NAND2_X1 U1564 ( .A1(n1937), .A2(G159), .ZN(n1439) );
  NAND2_X1 U1565 ( .A1(n1440), .A2(n1439), .ZN(n1444) );
  NAND2_X1 U1566 ( .A1(G143), .A2(n1921), .ZN(n1442) );
  NAND2_X1 U1567 ( .A1(G132), .A2(n1933), .ZN(n1441) );
  NAND2_X1 U1568 ( .A1(n1442), .A2(n1441), .ZN(n1443) );
  NOR2_X1 U1569 ( .A1(n1444), .A2(n1443), .ZN(n1452) );
  NOR2_X1 U1570 ( .A1(n1884), .A2(G33), .ZN(n1920) );
  NAND2_X1 U1571 ( .A1(n1927), .A2(G137), .ZN(n1445) );
  NAND2_X1 U1572 ( .A1(n1920), .A2(n1445), .ZN(n1450) );
  INV_X1 U1573 ( .A(n1446), .ZN(n1931) );
  NAND2_X1 U1574 ( .A1(G150), .A2(n1931), .ZN(n1448) );
  NAND2_X1 U1575 ( .A1(G50), .A2(n1928), .ZN(n1447) );
  NAND2_X1 U1576 ( .A1(n1448), .A2(n1447), .ZN(n1449) );
  NOR2_X1 U1577 ( .A1(n1450), .A2(n1449), .ZN(n1451) );
  NAND2_X1 U1578 ( .A1(n1452), .A2(n1451), .ZN(n1454) );
  NAND2_X1 U1579 ( .A1(G58), .A2(n1934), .ZN(n1453) );
  XNOR2_X1 U1580 ( .A(KEYINPUT97), .B(n1453), .ZN(n1859) );
  NOR2_X1 U1581 ( .A1(n1454), .A2(n1859), .ZN(n1455) );
  XOR2_X1 U1582 ( .A(KEYINPUT104), .B(n1455), .Z(n1456) );
  NAND2_X1 U1583 ( .A1(n1457), .A2(n1456), .ZN(n1458) );
  NOR2_X1 U1584 ( .A1(n1681), .A2(n1458), .ZN(n1459) );
  XNOR2_X1 U1585 ( .A(n1459), .B(KEYINPUT45), .ZN(n1461) );
  NOR2_X1 U1586 ( .A1(n1837), .A2(n1949), .ZN(n1460) );
  NOR2_X1 U1587 ( .A1(n1461), .A2(n1460), .ZN(n1464) );
  NOR2_X1 U1588 ( .A1(n1959), .A2(n1462), .ZN(n1463) );
  NOR2_X1 U1589 ( .A1(n1464), .A2(n1463), .ZN(n1465) );
  NAND2_X1 U1590 ( .A1(n1501), .A2(n1470), .ZN(n1482) );
  XNOR2_X1 U1591 ( .A(KEYINPUT72), .B(n1482), .ZN(n1471) );
  NAND2_X1 U1592 ( .A1(n1501), .A2(n1277), .ZN(n1472) );
  NAND2_X1 U1593 ( .A1(n1501), .A2(n1474), .ZN(n1475) );
  NAND2_X1 U1594 ( .A1(n1501), .A2(n1481), .ZN(n1477) );
  XNOR2_X2 U1595 ( .A(n1506), .B(n1503), .ZN(n1480) );
  NAND2_X1 U1596 ( .A1(n1501), .A2(n1479), .ZN(n1502) );
  XNOR2_X2 U1597 ( .A(n1480), .B(n1013), .ZN(n1793) );
  NAND2_X1 U1598 ( .A1(n1481), .A2(n1807), .ZN(n1483) );
  NAND2_X1 U1599 ( .A1(n1793), .A2(n1731), .ZN(n1486) );
  NAND2_X1 U1600 ( .A1(n1487), .A2(n1798), .ZN(n1489) );
  INV_X1 U1601 ( .A(KEYINPUT111), .ZN(n1488) );
  NAND2_X1 U1602 ( .A1(n1491), .A2(n1490), .ZN(n1493) );
  NAND2_X1 U1603 ( .A1(n1495), .A2(n1501), .ZN(n1496) );
  NOR2_X1 U1604 ( .A1(n1497), .A2(n1496), .ZN(n1498) );
  NOR2_X1 U1605 ( .A1(n1499), .A2(n1498), .ZN(n1510) );
  NAND2_X1 U1606 ( .A1(n1501), .A2(n1500), .ZN(n1505) );
  NAND2_X1 U1607 ( .A1(n1503), .A2(n1502), .ZN(n1504) );
  NAND2_X1 U1608 ( .A1(n1505), .A2(n1504), .ZN(n1784) );
  INV_X1 U1609 ( .A(n1506), .ZN(n1507) );
  NAND2_X1 U1610 ( .A1(n1784), .A2(n1507), .ZN(n1508) );
  XNOR2_X1 U1611 ( .A(n1508), .B(KEYINPUT112), .ZN(n1509) );
  XNOR2_X1 U1612 ( .A(n1510), .B(n1509), .ZN(n1511) );
  INV_X1 U1613 ( .A(n1681), .ZN(n1954) );
  NOR2_X1 U1614 ( .A1(n1949), .A2(G20), .ZN(n1534) );
  INV_X1 U1615 ( .A(n1534), .ZN(n1785) );
  NAND2_X1 U1616 ( .A1(n1884), .A2(n1785), .ZN(n1783) );
  NOR2_X1 U1617 ( .A1(n2002), .A2(n1740), .ZN(n1512) );
  XNOR2_X1 U1618 ( .A(n1512), .B(KEYINPUT24), .ZN(n1779) );
  XNOR2_X1 U1619 ( .A(G257), .B(G264), .ZN(n1513) );
  XNOR2_X1 U1620 ( .A(n1513), .B(G270), .ZN(n1514) );
  XNOR2_X1 U1621 ( .A(G250), .B(n1514), .ZN(n2058) );
  NAND2_X1 U1622 ( .A1(n1779), .A2(n2058), .ZN(n1516) );
  NAND2_X1 U1623 ( .A1(G87), .A2(n2002), .ZN(n1515) );
  NAND2_X1 U1624 ( .A1(n1516), .A2(n1515), .ZN(n1517) );
  NOR2_X1 U1625 ( .A1(n1783), .A2(n1517), .ZN(n1558) );
  NAND2_X1 U1626 ( .A1(G143), .A2(n1933), .ZN(n1519) );
  NAND2_X1 U1627 ( .A1(n1921), .A2(G159), .ZN(n1518) );
  NAND2_X1 U1628 ( .A1(n1519), .A2(n1518), .ZN(n1521) );
  NAND2_X1 U1629 ( .A1(G68), .A2(n1928), .ZN(n1846) );
  NAND2_X1 U1630 ( .A1(n1920), .A2(n1846), .ZN(n1520) );
  NOR2_X1 U1631 ( .A1(n1521), .A2(n1520), .ZN(n1532) );
  NAND2_X1 U1632 ( .A1(n1927), .A2(G150), .ZN(n1523) );
  NAND2_X1 U1633 ( .A1(n1931), .A2(G50), .ZN(n1522) );
  NAND2_X1 U1634 ( .A1(n1523), .A2(n1522), .ZN(n1530) );
  NAND2_X1 U1635 ( .A1(G137), .A2(n1922), .ZN(n1524) );
  XNOR2_X1 U1636 ( .A(n1524), .B(KEYINPUT115), .ZN(n1526) );
  INV_X1 U1637 ( .A(n1937), .ZN(n1564) );
  NOR2_X1 U1638 ( .A1(n1564), .A2(n1083), .ZN(n1525) );
  NOR2_X1 U1639 ( .A1(n1526), .A2(n1525), .ZN(n1528) );
  NAND2_X1 U1640 ( .A1(n1528), .A2(n1527), .ZN(n1529) );
  NOR2_X1 U1641 ( .A1(n1530), .A2(n1529), .ZN(n1531) );
  NAND2_X1 U1642 ( .A1(n1532), .A2(n1531), .ZN(n1536) );
  NAND2_X1 U1643 ( .A1(n1534), .A2(n1533), .ZN(n1535) );
  NAND2_X1 U1644 ( .A1(n1536), .A2(n1535), .ZN(n1555) );
  NOR2_X1 U1645 ( .A1(n1537), .A2(n1717), .ZN(n1553) );
  NAND2_X1 U1646 ( .A1(G97), .A2(n1934), .ZN(n1667) );
  NAND2_X1 U1647 ( .A1(n1922), .A2(G317), .ZN(n1538) );
  NAND2_X1 U1648 ( .A1(n1667), .A2(n1538), .ZN(n1540) );
  AND2_X1 U1649 ( .A1(G303), .A2(n1927), .ZN(n1539) );
  NOR2_X1 U1650 ( .A1(n1540), .A2(n1539), .ZN(n1547) );
  NAND2_X1 U1651 ( .A1(n1921), .A2(G294), .ZN(n1542) );
  NAND2_X1 U1652 ( .A1(n1937), .A2(G116), .ZN(n1541) );
  NAND2_X1 U1653 ( .A1(n1542), .A2(n1541), .ZN(n1545) );
  NAND2_X1 U1654 ( .A1(n1933), .A2(G311), .ZN(n1543) );
  XOR2_X1 U1655 ( .A(KEYINPUT54), .B(n1543), .Z(n1544) );
  NOR2_X1 U1656 ( .A1(n1545), .A2(n1544), .ZN(n1546) );
  NAND2_X1 U1657 ( .A1(n1547), .A2(n1546), .ZN(n1550) );
  NAND2_X1 U1658 ( .A1(G283), .A2(n1931), .ZN(n1548) );
  XOR2_X1 U1659 ( .A(KEYINPUT116), .B(n1548), .Z(n1549) );
  NOR2_X1 U1660 ( .A1(n1550), .A2(n1549), .ZN(n1551) );
  NAND2_X1 U1661 ( .A1(n1551), .A2(n1909), .ZN(n1552) );
  NOR2_X1 U1662 ( .A1(n1553), .A2(n1552), .ZN(n1554) );
  NOR2_X1 U1663 ( .A1(n1555), .A2(n1554), .ZN(n1556) );
  NAND2_X1 U1664 ( .A1(n1954), .A2(n1556), .ZN(n1557) );
  XOR2_X1 U1665 ( .A(n2019), .B(n1839), .Z(n1559) );
  NAND2_X1 U1666 ( .A1(n1559), .A2(n1681), .ZN(n1603) );
  NAND2_X1 U1667 ( .A1(G97), .A2(n1928), .ZN(n1640) );
  NAND2_X1 U1668 ( .A1(n1909), .A2(n1640), .ZN(n1571) );
  NAND2_X1 U1669 ( .A1(n1931), .A2(G116), .ZN(n1560) );
  XNOR2_X1 U1670 ( .A(n1560), .B(KEYINPUT21), .ZN(n1561) );
  XNOR2_X1 U1671 ( .A(KEYINPUT117), .B(n1561), .ZN(n1569) );
  NAND2_X1 U1672 ( .A1(n1933), .A2(G303), .ZN(n1563) );
  NAND2_X1 U1673 ( .A1(n1927), .A2(G294), .ZN(n1562) );
  NAND2_X1 U1674 ( .A1(n1563), .A2(n1562), .ZN(n1566) );
  NOR2_X1 U1675 ( .A1(n1717), .A2(n1564), .ZN(n1565) );
  NOR2_X1 U1676 ( .A1(n1566), .A2(n1565), .ZN(n1567) );
  XNOR2_X1 U1677 ( .A(KEYINPUT118), .B(n1567), .ZN(n1568) );
  NAND2_X1 U1678 ( .A1(n1569), .A2(n1568), .ZN(n1570) );
  NOR2_X1 U1679 ( .A1(n1571), .A2(n1570), .ZN(n1577) );
  NAND2_X1 U1680 ( .A1(G311), .A2(n1922), .ZN(n1573) );
  NAND2_X1 U1681 ( .A1(n1921), .A2(G283), .ZN(n1572) );
  NAND2_X1 U1682 ( .A1(n1573), .A2(n1572), .ZN(n1575) );
  NAND2_X1 U1683 ( .A1(n1934), .A2(G87), .ZN(n1574) );
  XOR2_X1 U1684 ( .A(KEYINPUT22), .B(n1574), .Z(n1766) );
  NOR2_X1 U1685 ( .A1(n1575), .A2(n1766), .ZN(n1576) );
  NAND2_X1 U1686 ( .A1(n1577), .A2(n1576), .ZN(n1578) );
  NAND2_X1 U1687 ( .A1(n1954), .A2(n1578), .ZN(n1580) );
  NOR2_X1 U1688 ( .A1(G77), .A2(n1899), .ZN(n1579) );
  NOR2_X1 U1689 ( .A1(n1580), .A2(n1579), .ZN(n1581) );
  XNOR2_X1 U1690 ( .A(n1581), .B(KEYINPUT119), .ZN(n1583) );
  NOR2_X1 U1691 ( .A1(n1949), .A2(n1839), .ZN(n1582) );
  NOR2_X1 U1692 ( .A1(n1583), .A2(n1582), .ZN(n1601) );
  NAND2_X1 U1693 ( .A1(n1927), .A2(G143), .ZN(n1584) );
  NAND2_X1 U1694 ( .A1(n1920), .A2(n1584), .ZN(n1593) );
  NAND2_X1 U1695 ( .A1(n1933), .A2(G137), .ZN(n1586) );
  NAND2_X1 U1696 ( .A1(G58), .A2(n1928), .ZN(n1585) );
  NAND2_X1 U1697 ( .A1(n1586), .A2(n1585), .ZN(n1590) );
  NAND2_X1 U1698 ( .A1(n1931), .A2(G159), .ZN(n1588) );
  NAND2_X1 U1699 ( .A1(n1937), .A2(G50), .ZN(n1587) );
  NAND2_X1 U1700 ( .A1(n1588), .A2(n1587), .ZN(n1589) );
  NOR2_X1 U1701 ( .A1(n1590), .A2(n1589), .ZN(n1591) );
  XOR2_X1 U1702 ( .A(KEYINPUT20), .B(n1591), .Z(n1592) );
  NOR2_X1 U1703 ( .A1(n1593), .A2(n1592), .ZN(n1599) );
  NAND2_X1 U1704 ( .A1(G68), .A2(n1934), .ZN(n1905) );
  NAND2_X1 U1705 ( .A1(G150), .A2(n1921), .ZN(n1594) );
  NAND2_X1 U1706 ( .A1(n1905), .A2(n1594), .ZN(n1597) );
  NAND2_X1 U1707 ( .A1(G132), .A2(n1922), .ZN(n1595) );
  XNOR2_X1 U1708 ( .A(n1595), .B(KEYINPUT19), .ZN(n1596) );
  NOR2_X1 U1709 ( .A1(n1597), .A2(n1596), .ZN(n1598) );
  NAND2_X1 U1710 ( .A1(n1599), .A2(n1598), .ZN(n1600) );
  NAND2_X1 U1711 ( .A1(n1601), .A2(n1600), .ZN(n1602) );
  NAND2_X1 U1712 ( .A1(n1603), .A2(n1602), .ZN(G384) );
  OR2_X1 U1713 ( .A1(n1605), .A2(n1604), .ZN(G355) );
  NAND2_X1 U1714 ( .A1(n1937), .A2(G303), .ZN(n1607) );
  NAND2_X1 U1715 ( .A1(n1934), .A2(G283), .ZN(n1606) );
  NAND2_X1 U1716 ( .A1(n1607), .A2(n1606), .ZN(n1620) );
  NAND2_X1 U1717 ( .A1(G317), .A2(n1921), .ZN(n1609) );
  NAND2_X1 U1718 ( .A1(G329), .A2(n1922), .ZN(n1608) );
  NAND2_X1 U1719 ( .A1(n1609), .A2(n1608), .ZN(n1611) );
  AND2_X1 U1720 ( .A1(n1928), .A2(G294), .ZN(n1610) );
  NOR2_X1 U1721 ( .A1(n1611), .A2(n1610), .ZN(n1618) );
  NAND2_X1 U1722 ( .A1(n1933), .A2(G326), .ZN(n1612) );
  NAND2_X1 U1723 ( .A1(n1909), .A2(n1612), .ZN(n1616) );
  NAND2_X1 U1724 ( .A1(G311), .A2(n1931), .ZN(n1614) );
  NAND2_X1 U1725 ( .A1(G322), .A2(n1927), .ZN(n1613) );
  NAND2_X1 U1726 ( .A1(n1614), .A2(n1613), .ZN(n1615) );
  NOR2_X1 U1727 ( .A1(n1616), .A2(n1615), .ZN(n1617) );
  NAND2_X1 U1728 ( .A1(n1618), .A2(n1617), .ZN(n1619) );
  NOR2_X1 U1729 ( .A1(n1620), .A2(n1619), .ZN(n1621) );
  NOR2_X1 U1730 ( .A1(n1681), .A2(n1621), .ZN(n1662) );
  NOR2_X1 U1731 ( .A1(n1622), .A2(n1785), .ZN(n1623) );
  XNOR2_X1 U1732 ( .A(n1623), .B(KEYINPUT62), .ZN(n1638) );
  NAND2_X1 U1733 ( .A1(n1080), .A2(n2002), .ZN(n1624) );
  XNOR2_X1 U1734 ( .A(n1624), .B(KEYINPUT60), .ZN(n1627) );
  INV_X1 U1735 ( .A(n1949), .ZN(n1625) );
  NAND2_X1 U1736 ( .A1(n1625), .A2(G355), .ZN(n1626) );
  NAND2_X1 U1737 ( .A1(n1627), .A2(n1626), .ZN(n1635) );
  XOR2_X1 U1738 ( .A(G77), .B(n2026), .Z(n1629) );
  XNOR2_X1 U1739 ( .A(n1629), .B(n1628), .ZN(n2061) );
  NAND2_X1 U1740 ( .A1(G45), .A2(n2061), .ZN(n1630) );
  NAND2_X1 U1741 ( .A1(n1779), .A2(n1630), .ZN(n1633) );
  NAND2_X1 U1742 ( .A1(n2052), .A2(G50), .ZN(n1631) );
  XNOR2_X1 U1743 ( .A(n1631), .B(KEYINPUT82), .ZN(n2015) );
  NOR2_X1 U1744 ( .A1(n2015), .A2(G45), .ZN(n1632) );
  NOR2_X1 U1745 ( .A1(n1633), .A2(n1632), .ZN(n1634) );
  NOR2_X1 U1746 ( .A1(n1635), .A2(n1634), .ZN(n1636) );
  NOR2_X1 U1747 ( .A1(n1783), .A2(n1636), .ZN(n1637) );
  NOR2_X1 U1748 ( .A1(n1638), .A2(n1637), .ZN(n1659) );
  NAND2_X1 U1749 ( .A1(n1922), .A2(G159), .ZN(n1646) );
  NAND2_X1 U1750 ( .A1(G77), .A2(n1931), .ZN(n1639) );
  NAND2_X1 U1751 ( .A1(n1640), .A2(n1639), .ZN(n1641) );
  XNOR2_X1 U1752 ( .A(KEYINPUT84), .B(n1641), .ZN(n1644) );
  NAND2_X1 U1753 ( .A1(G68), .A2(n1921), .ZN(n1642) );
  XNOR2_X1 U1754 ( .A(KEYINPUT83), .B(n1642), .ZN(n1643) );
  NOR2_X1 U1755 ( .A1(n1644), .A2(n1643), .ZN(n1645) );
  NAND2_X1 U1756 ( .A1(n1646), .A2(n1645), .ZN(n1647) );
  XNOR2_X1 U1757 ( .A(n1647), .B(KEYINPUT61), .ZN(n1653) );
  NAND2_X1 U1758 ( .A1(n1937), .A2(G87), .ZN(n1648) );
  XNOR2_X1 U1759 ( .A(n1648), .B(KEYINPUT85), .ZN(n1907) );
  NAND2_X1 U1760 ( .A1(G50), .A2(n1933), .ZN(n1649) );
  NAND2_X1 U1761 ( .A1(n1920), .A2(n1649), .ZN(n1650) );
  NOR2_X1 U1762 ( .A1(n1907), .A2(n1650), .ZN(n1651) );
  XNOR2_X1 U1763 ( .A(n1651), .B(KEYINPUT86), .ZN(n1652) );
  NAND2_X1 U1764 ( .A1(n1653), .A2(n1652), .ZN(n1656) );
  NOR2_X1 U1765 ( .A1(n1083), .A2(n1654), .ZN(n1655) );
  NOR2_X1 U1766 ( .A1(n1656), .A2(n1655), .ZN(n1657) );
  NAND2_X1 U1767 ( .A1(G107), .A2(n1934), .ZN(n1741) );
  NAND2_X1 U1768 ( .A1(n1657), .A2(n1741), .ZN(n1658) );
  NAND2_X1 U1769 ( .A1(n1659), .A2(n1658), .ZN(n1660) );
  XNOR2_X1 U1770 ( .A(KEYINPUT87), .B(n1660), .ZN(n1661) );
  NAND2_X1 U1771 ( .A1(n1662), .A2(n1661), .ZN(n1665) );
  XOR2_X1 U1772 ( .A(G330), .B(n1622), .Z(n1663) );
  NAND2_X1 U1773 ( .A1(n1663), .A2(n1681), .ZN(n1664) );
  NAND2_X1 U1774 ( .A1(n1665), .A2(n1664), .ZN(G396) );
  NAND2_X1 U1775 ( .A1(G159), .A2(n1933), .ZN(n1666) );
  NAND2_X1 U1776 ( .A1(n1667), .A2(n1666), .ZN(n1679) );
  NAND2_X1 U1777 ( .A1(G77), .A2(n1937), .ZN(n1853) );
  NAND2_X1 U1778 ( .A1(G150), .A2(n1922), .ZN(n1668) );
  NAND2_X1 U1779 ( .A1(n1853), .A2(n1668), .ZN(n1669) );
  NOR2_X1 U1780 ( .A1(n1670), .A2(n1669), .ZN(n1677) );
  NAND2_X1 U1781 ( .A1(G58), .A2(n1921), .ZN(n1671) );
  NAND2_X1 U1782 ( .A1(n1920), .A2(n1671), .ZN(n1675) );
  NAND2_X1 U1783 ( .A1(n1927), .A2(G50), .ZN(n1673) );
  NAND2_X1 U1784 ( .A1(n1931), .A2(G68), .ZN(n1672) );
  NAND2_X1 U1785 ( .A1(n1673), .A2(n1672), .ZN(n1674) );
  NOR2_X1 U1786 ( .A1(n1675), .A2(n1674), .ZN(n1676) );
  NAND2_X1 U1787 ( .A1(n1677), .A2(n1676), .ZN(n1678) );
  NOR2_X1 U1788 ( .A1(n1679), .A2(n1678), .ZN(n1680) );
  NOR2_X1 U1789 ( .A1(n1681), .A2(n1680), .ZN(n1685) );
  NOR2_X1 U1790 ( .A1(n1785), .A2(n1682), .ZN(n1683) );
  XNOR2_X1 U1791 ( .A(n1683), .B(KEYINPUT109), .ZN(n1684) );
  NAND2_X1 U1792 ( .A1(n1685), .A2(n1684), .ZN(n1727) );
  NAND2_X1 U1793 ( .A1(G317), .A2(n1927), .ZN(n1687) );
  NAND2_X1 U1794 ( .A1(n1931), .A2(G303), .ZN(n1686) );
  NAND2_X1 U1795 ( .A1(n1687), .A2(n1686), .ZN(n1699) );
  NAND2_X1 U1796 ( .A1(G326), .A2(n1922), .ZN(n1688) );
  XNOR2_X1 U1797 ( .A(n1688), .B(KEYINPUT105), .ZN(n1691) );
  NAND2_X1 U1798 ( .A1(G116), .A2(n1934), .ZN(n1689) );
  XNOR2_X1 U1799 ( .A(KEYINPUT25), .B(n1689), .ZN(n1690) );
  NOR2_X1 U1800 ( .A1(n1691), .A2(n1690), .ZN(n1697) );
  NAND2_X1 U1801 ( .A1(G283), .A2(n1928), .ZN(n1692) );
  NAND2_X1 U1802 ( .A1(n1909), .A2(n1692), .ZN(n1695) );
  NAND2_X1 U1803 ( .A1(n1921), .A2(G311), .ZN(n1693) );
  XOR2_X1 U1804 ( .A(KEYINPUT106), .B(n1693), .Z(n1694) );
  NOR2_X1 U1805 ( .A1(n1695), .A2(n1694), .ZN(n1696) );
  NAND2_X1 U1806 ( .A1(n1697), .A2(n1696), .ZN(n1698) );
  NOR2_X1 U1807 ( .A1(n1699), .A2(n1698), .ZN(n1704) );
  NAND2_X1 U1808 ( .A1(G322), .A2(n1933), .ZN(n1701) );
  NAND2_X1 U1809 ( .A1(n1937), .A2(G294), .ZN(n1700) );
  NAND2_X1 U1810 ( .A1(n1701), .A2(n1700), .ZN(n1702) );
  XOR2_X1 U1811 ( .A(KEYINPUT26), .B(n1702), .Z(n1703) );
  NAND2_X1 U1812 ( .A1(n1704), .A2(n1703), .ZN(n1725) );
  NOR2_X1 U1813 ( .A1(G116), .A2(n1705), .ZN(n2012) );
  NAND2_X1 U1814 ( .A1(n2012), .A2(n2026), .ZN(n1708) );
  NAND2_X1 U1815 ( .A1(G77), .A2(G68), .ZN(n1706) );
  NAND2_X1 U1816 ( .A1(G58), .A2(n1706), .ZN(n1707) );
  NOR2_X1 U1817 ( .A1(n1708), .A2(n1707), .ZN(n1709) );
  NOR2_X1 U1818 ( .A1(G45), .A2(n1709), .ZN(n1710) );
  XNOR2_X1 U1819 ( .A(n1710), .B(KEYINPUT23), .ZN(n1715) );
  XOR2_X1 U1820 ( .A(KEYINPUT107), .B(G226), .Z(n1712) );
  XNOR2_X1 U1821 ( .A(G244), .B(G232), .ZN(n1711) );
  XNOR2_X1 U1822 ( .A(n1712), .B(n1711), .ZN(n1713) );
  XOR2_X1 U1823 ( .A(G238), .B(n1713), .Z(n2059) );
  NAND2_X1 U1824 ( .A1(n2059), .A2(G45), .ZN(n1714) );
  NAND2_X1 U1825 ( .A1(n1715), .A2(n1714), .ZN(n1716) );
  NAND2_X1 U1826 ( .A1(n1716), .A2(n1779), .ZN(n1719) );
  NAND2_X1 U1827 ( .A1(n2002), .A2(n1717), .ZN(n1718) );
  NAND2_X1 U1828 ( .A1(n1719), .A2(n1718), .ZN(n1721) );
  NOR2_X1 U1829 ( .A1(n2012), .A2(n1949), .ZN(n1720) );
  NOR2_X1 U1830 ( .A1(n1721), .A2(n1720), .ZN(n1722) );
  NOR2_X1 U1831 ( .A1(n1783), .A2(n1722), .ZN(n1723) );
  XOR2_X1 U1832 ( .A(KEYINPUT108), .B(n1723), .Z(n1724) );
  NAND2_X1 U1833 ( .A1(n1725), .A2(n1724), .ZN(n1726) );
  NOR2_X1 U1834 ( .A1(n1727), .A2(n1726), .ZN(n1729) );
  INV_X1 U1835 ( .A(n1731), .ZN(n1794) );
  NOR2_X1 U1836 ( .A1(n1736), .A2(n1794), .ZN(n1728) );
  NOR2_X1 U1837 ( .A1(n1729), .A2(n1728), .ZN(n1734) );
  NOR2_X1 U1838 ( .A1(n2014), .A2(n1731), .ZN(n1732) );
  NAND2_X1 U1839 ( .A1(n1730), .A2(n1732), .ZN(n1733) );
  NAND2_X1 U1840 ( .A1(n1734), .A2(n1733), .ZN(G393) );
  INV_X1 U1841 ( .A(n1793), .ZN(n1735) );
  NOR2_X1 U1842 ( .A1(n1736), .A2(n1735), .ZN(n1792) );
  NAND2_X1 U1843 ( .A1(G322), .A2(n1922), .ZN(n1738) );
  NAND2_X1 U1844 ( .A1(G311), .A2(n1927), .ZN(n1737) );
  NAND2_X1 U1845 ( .A1(n1738), .A2(n1737), .ZN(n1739) );
  NOR2_X1 U1846 ( .A1(n1740), .A2(n1739), .ZN(n1748) );
  NAND2_X1 U1847 ( .A1(G303), .A2(n1921), .ZN(n1742) );
  NAND2_X1 U1848 ( .A1(n1742), .A2(n1741), .ZN(n1746) );
  NAND2_X1 U1849 ( .A1(G294), .A2(n1931), .ZN(n1744) );
  NAND2_X1 U1850 ( .A1(G116), .A2(n1928), .ZN(n1743) );
  NAND2_X1 U1851 ( .A1(n1744), .A2(n1743), .ZN(n1745) );
  NOR2_X1 U1852 ( .A1(n1746), .A2(n1745), .ZN(n1747) );
  NAND2_X1 U1853 ( .A1(n1748), .A2(n1747), .ZN(n1749) );
  XNOR2_X1 U1854 ( .A(KEYINPUT58), .B(n1749), .ZN(n1755) );
  NAND2_X1 U1855 ( .A1(n1933), .A2(G317), .ZN(n1750) );
  XOR2_X1 U1856 ( .A(KEYINPUT79), .B(n1750), .Z(n1752) );
  NAND2_X1 U1857 ( .A1(G283), .A2(n1937), .ZN(n1751) );
  NAND2_X1 U1858 ( .A1(n1752), .A2(n1751), .ZN(n1753) );
  XOR2_X1 U1859 ( .A(KEYINPUT59), .B(n1753), .Z(n1754) );
  NOR2_X1 U1860 ( .A1(n1755), .A2(n1754), .ZN(n1773) );
  NAND2_X1 U1861 ( .A1(G143), .A2(n1922), .ZN(n1757) );
  NAND2_X1 U1862 ( .A1(n1921), .A2(G50), .ZN(n1756) );
  NAND2_X1 U1863 ( .A1(n1757), .A2(n1756), .ZN(n1760) );
  NAND2_X1 U1864 ( .A1(G58), .A2(n1931), .ZN(n1758) );
  NAND2_X1 U1865 ( .A1(n1861), .A2(n1758), .ZN(n1759) );
  NOR2_X1 U1866 ( .A1(n1760), .A2(n1759), .ZN(n1768) );
  NAND2_X1 U1867 ( .A1(G150), .A2(n1933), .ZN(n1761) );
  XNOR2_X1 U1868 ( .A(n1761), .B(KEYINPUT56), .ZN(n1763) );
  NAND2_X1 U1869 ( .A1(n1937), .A2(G68), .ZN(n1762) );
  NAND2_X1 U1870 ( .A1(n1763), .A2(n1762), .ZN(n1764) );
  XOR2_X1 U1871 ( .A(KEYINPUT57), .B(n1764), .Z(n1765) );
  NOR2_X1 U1872 ( .A1(n1766), .A2(n1765), .ZN(n1767) );
  NAND2_X1 U1873 ( .A1(n1768), .A2(n1767), .ZN(n1771) );
  NAND2_X1 U1874 ( .A1(G77), .A2(n1928), .ZN(n1908) );
  NAND2_X1 U1875 ( .A1(G159), .A2(n1927), .ZN(n1769) );
  NAND2_X1 U1876 ( .A1(n1908), .A2(n1769), .ZN(n1770) );
  NOR2_X1 U1877 ( .A1(n1771), .A2(n1770), .ZN(n1772) );
  NOR2_X1 U1878 ( .A1(n1773), .A2(n1772), .ZN(n1774) );
  XNOR2_X1 U1879 ( .A(n1774), .B(KEYINPUT80), .ZN(n1775) );
  NOR2_X1 U1880 ( .A1(n1884), .A2(n1775), .ZN(n1790) );
  XNOR2_X1 U1881 ( .A(n1080), .B(KEYINPUT51), .ZN(n1776) );
  XNOR2_X1 U1882 ( .A(n2023), .B(n1776), .ZN(n1777) );
  XOR2_X1 U1883 ( .A(n1778), .B(n1777), .Z(n2060) );
  NAND2_X1 U1884 ( .A1(n1779), .A2(n2060), .ZN(n1781) );
  NAND2_X1 U1885 ( .A1(G97), .A2(n2002), .ZN(n1780) );
  NAND2_X1 U1886 ( .A1(n1781), .A2(n1780), .ZN(n1782) );
  NOR2_X1 U1887 ( .A1(n1783), .A2(n1782), .ZN(n1787) );
  NOR2_X1 U1888 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  NOR2_X1 U1889 ( .A1(n1787), .A2(n1786), .ZN(n1788) );
  NAND2_X1 U1890 ( .A1(n1954), .A2(n1788), .ZN(n1789) );
  NOR2_X1 U1891 ( .A1(n1790), .A2(n1789), .ZN(n1791) );
  NOR2_X1 U1892 ( .A1(n1792), .A2(n1791), .ZN(n1800) );
  NOR2_X1 U1893 ( .A1(n2019), .A2(n1794), .ZN(n1795) );
  NOR2_X1 U1894 ( .A1(n1793), .A2(n1795), .ZN(n1796) );
  NOR2_X1 U1895 ( .A1(n2014), .A2(n1796), .ZN(n1797) );
  NAND2_X1 U1896 ( .A1(n1798), .A2(n1797), .ZN(n1799) );
  NAND2_X1 U1897 ( .A1(n1800), .A2(n1799), .ZN(G390) );
  NAND2_X1 U1898 ( .A1(n1801), .A2(n1837), .ZN(n1802) );
  NAND2_X1 U1899 ( .A1(n1803), .A2(n1837), .ZN(n1804) );
  NAND2_X1 U1900 ( .A1(n1805), .A2(n1804), .ZN(n1806) );
  AND2_X1 U1901 ( .A1(n1807), .A2(n1806), .ZN(n1832) );
  NAND2_X1 U1902 ( .A1(n1809), .A2(n1834), .ZN(n1811) );
  NAND2_X1 U1903 ( .A1(n1811), .A2(n1810), .ZN(n1814) );
  NAND2_X1 U1904 ( .A1(n1812), .A2(n1834), .ZN(n1813) );
  NAND2_X1 U1905 ( .A1(n1814), .A2(n1813), .ZN(n1815) );
  XNOR2_X1 U1906 ( .A(n1819), .B(n1818), .ZN(n1960) );
  NAND2_X1 U1907 ( .A1(n1960), .A2(n1897), .ZN(n1821) );
  XOR2_X1 U1908 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n1820) );
  XNOR2_X1 U1909 ( .A(n1821), .B(n1820), .ZN(n1824) );
  NOR2_X1 U1910 ( .A1(n1822), .A2(n1068), .ZN(n1823) );
  NAND2_X1 U1911 ( .A1(n1825), .A2(n1834), .ZN(n1828) );
  INV_X1 U1912 ( .A(n1826), .ZN(n1827) );
  NAND2_X1 U1913 ( .A1(n1828), .A2(n1827), .ZN(n1831) );
  NAND2_X1 U1914 ( .A1(n1829), .A2(n1834), .ZN(n1830) );
  NAND2_X1 U1915 ( .A1(n1831), .A2(n1830), .ZN(n1891) );
  AND2_X1 U1916 ( .A1(n1950), .A2(n1832), .ZN(n1836) );
  NOR2_X1 U1917 ( .A1(n1834), .A2(n1833), .ZN(n1835) );
  NOR2_X1 U1918 ( .A1(n1836), .A2(n1835), .ZN(n2039) );
  NAND2_X1 U1919 ( .A1(n1837), .A2(n1950), .ZN(n1841) );
  NAND2_X1 U1920 ( .A1(n1838), .A2(n1839), .ZN(n1840) );
  NOR2_X1 U1921 ( .A1(n1841), .A2(n1840), .ZN(n2037) );
  NAND2_X1 U1922 ( .A1(G330), .A2(n2037), .ZN(n1842) );
  NAND2_X1 U1923 ( .A1(n2039), .A2(n1842), .ZN(n1843) );
  XOR2_X1 U1924 ( .A(n1891), .B(n1843), .Z(n1844) );
  NAND2_X1 U1925 ( .A1(n1089), .A2(n1090), .ZN(n1896) );
  NAND2_X1 U1926 ( .A1(G87), .A2(n1931), .ZN(n1845) );
  NAND2_X1 U1927 ( .A1(n1846), .A2(n1845), .ZN(n1849) );
  NAND2_X1 U1928 ( .A1(G107), .A2(n1927), .ZN(n1847) );
  XOR2_X1 U1929 ( .A(KEYINPUT42), .B(n1847), .Z(n1848) );
  NOR2_X1 U1930 ( .A1(n1849), .A2(n1848), .ZN(n1857) );
  NAND2_X1 U1931 ( .A1(n1933), .A2(G116), .ZN(n1851) );
  NAND2_X1 U1932 ( .A1(n1921), .A2(G97), .ZN(n1850) );
  NAND2_X1 U1933 ( .A1(n1851), .A2(n1850), .ZN(n1855) );
  NAND2_X1 U1934 ( .A1(G283), .A2(n1922), .ZN(n1852) );
  NAND2_X1 U1935 ( .A1(n1853), .A2(n1852), .ZN(n1854) );
  NOR2_X1 U1936 ( .A1(n1855), .A2(n1854), .ZN(n1856) );
  NAND2_X1 U1937 ( .A1(n1857), .A2(n1856), .ZN(n1858) );
  NOR2_X1 U1938 ( .A1(n1859), .A2(n1858), .ZN(n1860) );
  NOR2_X1 U1939 ( .A1(n1861), .A2(n1860), .ZN(n1883) );
  NAND2_X1 U1940 ( .A1(n1921), .A2(G132), .ZN(n1862) );
  XNOR2_X1 U1941 ( .A(n1862), .B(KEYINPUT94), .ZN(n1864) );
  NAND2_X1 U1942 ( .A1(n1934), .A2(G159), .ZN(n1863) );
  NAND2_X1 U1943 ( .A1(n1864), .A2(n1863), .ZN(n1866) );
  XOR2_X1 U1944 ( .A(KEYINPUT44), .B(KEYINPUT95), .Z(n1865) );
  XNOR2_X1 U1945 ( .A(n1866), .B(n1865), .ZN(n1880) );
  NAND2_X1 U1946 ( .A1(G125), .A2(n1933), .ZN(n1868) );
  NAND2_X1 U1947 ( .A1(G143), .A2(n1937), .ZN(n1867) );
  NAND2_X1 U1948 ( .A1(n1868), .A2(n1867), .ZN(n1872) );
  NAND2_X1 U1949 ( .A1(G124), .A2(n1922), .ZN(n1870) );
  NAND2_X1 U1950 ( .A1(G128), .A2(n1927), .ZN(n1869) );
  NAND2_X1 U1951 ( .A1(n1870), .A2(n1869), .ZN(n1871) );
  NOR2_X1 U1952 ( .A1(n1872), .A2(n1871), .ZN(n1878) );
  NAND2_X1 U1953 ( .A1(n1928), .A2(G150), .ZN(n1873) );
  XOR2_X1 U1954 ( .A(KEYINPUT96), .B(n1873), .Z(n1876) );
  NAND2_X1 U1955 ( .A1(G137), .A2(n1931), .ZN(n1874) );
  XNOR2_X1 U1956 ( .A(KEYINPUT43), .B(n1874), .ZN(n1875) );
  NOR2_X1 U1957 ( .A1(n1876), .A2(n1875), .ZN(n1877) );
  NAND2_X1 U1958 ( .A1(n1878), .A2(n1877), .ZN(n1879) );
  NOR2_X1 U1959 ( .A1(n1880), .A2(n1879), .ZN(n1881) );
  NOR2_X1 U1960 ( .A1(G33), .A2(n1881), .ZN(n1882) );
  NOR2_X1 U1961 ( .A1(n1883), .A2(n1882), .ZN(n1885) );
  NOR2_X1 U1962 ( .A1(G41), .A2(n1884), .ZN(n1886) );
  NAND2_X1 U1963 ( .A1(n1885), .A2(n1886), .ZN(n1889) );
  NOR2_X1 U1964 ( .A1(G50), .A2(n1886), .ZN(n1887) );
  NAND2_X1 U1965 ( .A1(n1887), .A2(n1949), .ZN(n1888) );
  NAND2_X1 U1966 ( .A1(n1889), .A2(n1888), .ZN(n1890) );
  XNOR2_X1 U1967 ( .A(n1890), .B(KEYINPUT98), .ZN(n1893) );
  NOR2_X1 U1968 ( .A1(n1891), .A2(n1949), .ZN(n1892) );
  NOR2_X1 U1969 ( .A1(n1893), .A2(n1892), .ZN(n1894) );
  NAND2_X1 U1970 ( .A1(n1894), .A2(n1954), .ZN(n1895) );
  NAND2_X1 U1971 ( .A1(n1896), .A2(n1895), .ZN(G375) );
  NOR2_X1 U1972 ( .A1(n2014), .A2(n1898), .ZN(n1958) );
  NOR2_X1 U1973 ( .A1(G58), .A2(n1899), .ZN(n1956) );
  NAND2_X1 U1974 ( .A1(n1922), .A2(G294), .ZN(n1901) );
  NAND2_X1 U1975 ( .A1(n1931), .A2(G97), .ZN(n1900) );
  NAND2_X1 U1976 ( .A1(n1901), .A2(n1900), .ZN(n1903) );
  XOR2_X1 U1977 ( .A(KEYINPUT48), .B(KEYINPUT102), .Z(n1902) );
  XNOR2_X1 U1978 ( .A(n1903), .B(n1902), .ZN(n1919) );
  NAND2_X1 U1979 ( .A1(G107), .A2(n1921), .ZN(n1904) );
  NAND2_X1 U1980 ( .A1(n1905), .A2(n1904), .ZN(n1906) );
  NOR2_X1 U1981 ( .A1(n1907), .A2(n1906), .ZN(n1914) );
  NAND2_X1 U1982 ( .A1(n1909), .A2(n1908), .ZN(n1912) );
  NAND2_X1 U1983 ( .A1(G283), .A2(n1933), .ZN(n1910) );
  XNOR2_X1 U1984 ( .A(KEYINPUT101), .B(n1910), .ZN(n1911) );
  NOR2_X1 U1985 ( .A1(n1912), .A2(n1911), .ZN(n1913) );
  NAND2_X1 U1986 ( .A1(n1914), .A2(n1913), .ZN(n1917) );
  NAND2_X1 U1987 ( .A1(G116), .A2(n1927), .ZN(n1915) );
  XNOR2_X1 U1988 ( .A(KEYINPUT47), .B(n1915), .ZN(n1916) );
  NOR2_X1 U1989 ( .A1(n1917), .A2(n1916), .ZN(n1918) );
  NAND2_X1 U1990 ( .A1(n1919), .A2(n1918), .ZN(n1948) );
  INV_X1 U1991 ( .A(n1920), .ZN(n1926) );
  NAND2_X1 U1992 ( .A1(G137), .A2(n1921), .ZN(n1924) );
  NAND2_X1 U1993 ( .A1(G125), .A2(n1922), .ZN(n1923) );
  NAND2_X1 U1994 ( .A1(n1924), .A2(n1923), .ZN(n1925) );
  NOR2_X1 U1995 ( .A1(n1926), .A2(n1925), .ZN(n1946) );
  NAND2_X1 U1996 ( .A1(n1927), .A2(G132), .ZN(n1930) );
  NAND2_X1 U1997 ( .A1(G159), .A2(n1928), .ZN(n1929) );
  NAND2_X1 U1998 ( .A1(n1930), .A2(n1929), .ZN(n1944) );
  NAND2_X1 U1999 ( .A1(G143), .A2(n1931), .ZN(n1932) );
  XNOR2_X1 U2000 ( .A(n1932), .B(KEYINPUT100), .ZN(n1942) );
  NAND2_X1 U2001 ( .A1(G128), .A2(n1933), .ZN(n1936) );
  NAND2_X1 U2002 ( .A1(n1934), .A2(G50), .ZN(n1935) );
  NAND2_X1 U2003 ( .A1(n1936), .A2(n1935), .ZN(n1940) );
  NAND2_X1 U2004 ( .A1(G150), .A2(n1937), .ZN(n1938) );
  XNOR2_X1 U2005 ( .A(KEYINPUT99), .B(n1938), .ZN(n1939) );
  NOR2_X1 U2006 ( .A1(n1940), .A2(n1939), .ZN(n1941) );
  NAND2_X1 U2007 ( .A1(n1942), .A2(n1941), .ZN(n1943) );
  NOR2_X1 U2008 ( .A1(n1944), .A2(n1943), .ZN(n1945) );
  NAND2_X1 U2009 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
  NAND2_X1 U2010 ( .A1(n1948), .A2(n1947), .ZN(n1952) );
  NOR2_X1 U2011 ( .A1(n1950), .A2(n1949), .ZN(n1951) );
  NOR2_X1 U2012 ( .A1(n1952), .A2(n1951), .ZN(n1953) );
  NAND2_X1 U2013 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  NOR2_X1 U2014 ( .A1(n1956), .A2(n1955), .ZN(n1957) );
  NOR2_X1 U2015 ( .A1(n1958), .A2(n1957), .ZN(n1962) );
  NAND2_X1 U2016 ( .A1(n1960), .A2(n1068), .ZN(n1961) );
  NAND2_X1 U2017 ( .A1(n1962), .A2(n1961), .ZN(G378) );
  XNOR2_X1 U2018 ( .A(G381), .B(G387), .ZN(n1966) );
  XNOR2_X1 U2019 ( .A(G393), .B(G390), .ZN(n1964) );
  XNOR2_X1 U2020 ( .A(n1966), .B(n1965), .ZN(n2062) );
  XNOR2_X1 U2021 ( .A(n2062), .B(KEYINPUT120), .ZN(n1972) );
  INV_X1 U2022 ( .A(G213), .ZN(n1980) );
  NOR2_X1 U2023 ( .A1(G343), .A2(n1980), .ZN(n1967) );
  NOR2_X1 U2024 ( .A1(n2063), .A2(n1967), .ZN(n1970) );
  NAND2_X1 U2025 ( .A1(n1967), .A2(G2897), .ZN(n1968) );
  XNOR2_X1 U2026 ( .A(n1968), .B(KEYINPUT63), .ZN(n1969) );
  XNOR2_X1 U2027 ( .A(n1972), .B(n1971), .ZN(G405) );
  NOR2_X1 U2028 ( .A1(G393), .A2(G390), .ZN(n1977) );
  OR2_X1 U2029 ( .A1(G375), .A2(G378), .ZN(n1978) );
  NOR2_X1 U2030 ( .A1(G387), .A2(G381), .ZN(n1974) );
  NOR2_X1 U2031 ( .A1(G384), .A2(G396), .ZN(n1973) );
  NAND2_X1 U2032 ( .A1(n1974), .A2(n1973), .ZN(n1975) );
  NOR2_X1 U2033 ( .A1(n1978), .A2(n1975), .ZN(n1976) );
  NAND2_X1 U2034 ( .A1(n1977), .A2(n1976), .ZN(G407) );
  NOR2_X1 U2035 ( .A1(G343), .A2(n1978), .ZN(n1979) );
  NOR2_X1 U2036 ( .A1(n1980), .A2(n1979), .ZN(n1981) );
  NAND2_X1 U2037 ( .A1(n1981), .A2(G407), .ZN(G409) );
  NAND2_X1 U2038 ( .A1(G97), .A2(G257), .ZN(n1999) );
  NAND2_X1 U2039 ( .A1(G270), .A2(G116), .ZN(n1983) );
  NAND2_X1 U2040 ( .A1(G250), .A2(G87), .ZN(n1982) );
  NAND2_X1 U2041 ( .A1(n1983), .A2(n1982), .ZN(n1997) );
  NAND2_X1 U2042 ( .A1(G264), .A2(G107), .ZN(n1984) );
  XNOR2_X1 U2043 ( .A(n1984), .B(KEYINPUT50), .ZN(n1995) );
  NAND2_X1 U2044 ( .A1(G226), .A2(G50), .ZN(n1986) );
  NAND2_X1 U2045 ( .A1(G58), .A2(G232), .ZN(n1985) );
  NAND2_X1 U2046 ( .A1(n1986), .A2(n1985), .ZN(n1987) );
  XNOR2_X1 U2047 ( .A(n1987), .B(KEYINPUT121), .ZN(n1989) );
  NAND2_X1 U2048 ( .A1(G77), .A2(G244), .ZN(n1988) );
  NAND2_X1 U2049 ( .A1(n1989), .A2(n1988), .ZN(n1992) );
  NAND2_X1 U2050 ( .A1(G238), .A2(G68), .ZN(n1990) );
  XOR2_X1 U2051 ( .A(KEYINPUT122), .B(n1990), .Z(n1991) );
  NOR2_X1 U2052 ( .A1(n1992), .A2(n1991), .ZN(n1993) );
  XOR2_X1 U2053 ( .A(KEYINPUT49), .B(n1993), .Z(n1994) );
  NAND2_X1 U2054 ( .A1(n1995), .A2(n1994), .ZN(n1996) );
  NOR2_X1 U2055 ( .A1(n1997), .A2(n1996), .ZN(n1998) );
  NAND2_X1 U2056 ( .A1(n1999), .A2(n1998), .ZN(n2001) );
  INV_X1 U2057 ( .A(n1405), .ZN(n2000) );
  NAND2_X1 U2058 ( .A1(n2001), .A2(n2000), .ZN(n2006) );
  NOR2_X1 U2059 ( .A1(G257), .A2(G264), .ZN(n2003) );
  NOR2_X1 U2060 ( .A1(n2003), .A2(n2002), .ZN(n2004) );
  NAND2_X1 U2061 ( .A1(G250), .A2(n2004), .ZN(n2005) );
  NAND2_X1 U2062 ( .A1(n2006), .A2(n2005), .ZN(n2009) );
  NAND2_X1 U2063 ( .A1(G20), .A2(n2007), .ZN(n2043) );
  NOR2_X1 U2064 ( .A1(n2015), .A2(n2043), .ZN(n2008) );
  NOR2_X1 U2065 ( .A1(n2009), .A2(n2008), .ZN(G361) );
  AND2_X1 U2066 ( .A1(n2010), .A2(n2035), .ZN(G372) );
  NAND2_X1 U2067 ( .A1(n2011), .A2(n1506), .ZN(G399) );
  NAND2_X1 U2068 ( .A1(n2012), .A2(G1), .ZN(n2013) );
  NAND2_X1 U2069 ( .A1(n2014), .A2(n2013), .ZN(n2018) );
  NAND2_X1 U2070 ( .A1(n2016), .A2(n2015), .ZN(n2017) );
  NAND2_X1 U2071 ( .A1(n2018), .A2(n2017), .ZN(n2022) );
  NAND2_X1 U2072 ( .A1(n2020), .A2(n2019), .ZN(n2021) );
  NAND2_X1 U2073 ( .A1(n2022), .A2(n2021), .ZN(G364) );
  NOR2_X1 U2074 ( .A1(n2023), .A2(n2043), .ZN(n2024) );
  NAND2_X1 U2075 ( .A1(G116), .A2(n2024), .ZN(n2025) );
  XNOR2_X1 U2076 ( .A(KEYINPUT126), .B(n2025), .ZN(n2050) );
  NOR2_X1 U2077 ( .A1(G77), .A2(n2026), .ZN(n2027) );
  XNOR2_X1 U2078 ( .A(n2027), .B(KEYINPUT124), .ZN(n2030) );
  NAND2_X1 U2079 ( .A1(G58), .A2(G50), .ZN(n2028) );
  XOR2_X1 U2080 ( .A(G68), .B(n2028), .Z(n2029) );
  NOR2_X1 U2081 ( .A1(n2030), .A2(n2029), .ZN(n2032) );
  NAND2_X1 U2082 ( .A1(G1), .A2(n2031), .ZN(n2045) );
  NOR2_X1 U2083 ( .A1(n2032), .A2(n2045), .ZN(n2033) );
  XNOR2_X1 U2084 ( .A(n2033), .B(KEYINPUT125), .ZN(n2048) );
  NAND2_X1 U2085 ( .A1(n1838), .A2(n2035), .ZN(n2036) );
  XNOR2_X1 U2086 ( .A(n2037), .B(n2036), .ZN(n2038) );
  NAND2_X1 U2087 ( .A1(n2038), .A2(G330), .ZN(n2041) );
  XOR2_X1 U2088 ( .A(n2039), .B(KEYINPUT123), .Z(n2040) );
  XNOR2_X1 U2089 ( .A(n2041), .B(n2040), .ZN(n2042) );
  XNOR2_X1 U2090 ( .A(n2034), .B(n2042), .ZN(n2044) );
  NAND2_X1 U2091 ( .A1(n2044), .A2(n2043), .ZN(n2046) );
  NAND2_X1 U2092 ( .A1(n2046), .A2(n2045), .ZN(n2047) );
  NAND2_X1 U2093 ( .A1(n2048), .A2(n2047), .ZN(n2049) );
  NAND2_X1 U2094 ( .A1(n2050), .A2(n2049), .ZN(G367) );
  OR2_X1 U2095 ( .A1(G77), .A2(G50), .ZN(n2051) );
  NOR2_X1 U2096 ( .A1(n2052), .A2(n2051), .ZN(G353) );
  XNOR2_X1 U2097 ( .A(KEYINPUT127), .B(n2054), .ZN(n2057) );
  INV_X1 U2098 ( .A(n2055), .ZN(n2056) );
  NAND2_X1 U2099 ( .A1(n2057), .A2(n2056), .ZN(G369) );
  XOR2_X1 U2100 ( .A(n2059), .B(n2058), .Z(G358) );
  XNOR2_X1 U2101 ( .A(n2061), .B(n2060), .ZN(G351) );
  XNOR2_X1 U2102 ( .A(n2063), .B(n2062), .ZN(G402) );
endmodule

