//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G131), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT69), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G237), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G953), .ZN(new_n197));
  AND4_X1   g011(.A1(G143), .A2(new_n196), .A3(G214), .A4(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(G953), .B1(new_n193), .B2(new_n195), .ZN(new_n199));
  AOI21_X1  g013(.A(G143), .B1(new_n199), .B2(G214), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n191), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n194), .A2(G237), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n192), .A2(KEYINPUT69), .ZN(new_n205));
  OAI211_X1 g019(.A(G214), .B(new_n197), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(G143), .A3(G214), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n190), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(new_n202), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  XOR2_X1   g027(.A(G125), .B(G140), .Z(new_n214));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(G146), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n190), .B1(new_n208), .B2(new_n209), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n203), .A2(new_n211), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G113), .B(G122), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT18), .B(G131), .C1(new_n198), .C2(new_n200), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n214), .A2(KEYINPUT77), .A3(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n230));
  XNOR2_X1  g044(.A(G125), .B(G140), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n217), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n229), .A2(new_n232), .B1(new_n217), .B2(new_n231), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT18), .A2(G131), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n208), .A2(new_n209), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n224), .A2(new_n227), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT92), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n198), .A2(new_n200), .A3(new_n191), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n222), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n201), .A2(KEYINPUT92), .A3(new_n210), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n214), .B(KEYINPUT19), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n219), .B1(new_n242), .B2(G146), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n227), .B1(new_n245), .B2(new_n236), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n187), .B(new_n188), .C1(new_n237), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n224), .A2(new_n227), .A3(new_n236), .ZN(new_n248));
  INV_X1    g062(.A(new_n236), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n201), .A2(new_n210), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n243), .B1(new_n250), .B2(new_n238), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n251), .B2(new_n241), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n252), .B2(new_n227), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n187), .B1(new_n253), .B2(new_n188), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT94), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n247), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n253), .A2(KEYINPUT94), .A3(new_n187), .A4(new_n188), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n224), .A2(new_n236), .ZN(new_n259));
  INV_X1    g073(.A(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(G902), .B1(new_n261), .B2(new_n248), .ZN(new_n262));
  INV_X1    g076(.A(G475), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n207), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n207), .A2(G128), .ZN(new_n268));
  OR3_X1    g082(.A1(new_n267), .A2(new_n268), .A3(G134), .ZN(new_n269));
  XNOR2_X1  g083(.A(G116), .B(G122), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT13), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n266), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n276), .A2(KEYINPUT95), .B1(KEYINPUT13), .B2(new_n267), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(KEYINPUT95), .B2(new_n276), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n274), .B1(new_n278), .B2(G134), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT14), .A3(G122), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G107), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n270), .ZN(new_n284));
  OAI21_X1  g098(.A(G134), .B1(new_n267), .B2(new_n268), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n272), .B(new_n284), .C1(new_n269), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT9), .B(G234), .ZN(new_n288));
  INV_X1    g102(.A(G217), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(G953), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n287), .B(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G478), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(KEYINPUT15), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n291), .B(new_n292), .C1(KEYINPUT15), .C2(new_n294), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G952), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(G234), .A2(G237), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT21), .B(G898), .Z(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(G902), .A3(G953), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT96), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n258), .A2(new_n265), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G128), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n217), .A2(G143), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n207), .A2(G146), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G143), .B(G146), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT67), .A3(new_n313), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(G128), .B1(new_n314), .B2(new_n315), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n207), .A2(KEYINPUT1), .A3(G146), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n212), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT0), .A2(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT0), .B(G128), .Z(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(G125), .C1(new_n319), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n197), .A2(G224), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n271), .A3(G104), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n226), .A2(G107), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n226), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n271), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(KEYINPUT2), .A2(G113), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT2), .A2(G113), .ZN(new_n345));
  AND2_X1   g159(.A1(G116), .A2(G119), .ZN(new_n346));
  NOR2_X1   g160(.A1(G116), .A2(G119), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT5), .B1(new_n346), .B2(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n352));
  INV_X1    g166(.A(G119), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G116), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT87), .A4(G116), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n356), .A3(G113), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G101), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(KEYINPUT81), .A3(G101), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n344), .A2(new_n345), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n346), .A2(new_n347), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n348), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n371), .A3(G101), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n334), .B(new_n359), .C1(new_n366), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT6), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n359), .B1(new_n366), .B2(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(new_n334), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n380), .A3(new_n377), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n333), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n334), .B(KEYINPUT8), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n351), .B(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n356), .A2(G113), .A3(new_n357), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n349), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n358), .A2(new_n348), .B1(new_n340), .B2(new_n343), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n332), .A2(KEYINPUT7), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n326), .B(new_n330), .C1(KEYINPUT90), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n330), .B2(KEYINPUT90), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n331), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n374), .A2(new_n391), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n292), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n311), .B1(new_n384), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n396), .A2(new_n292), .ZN(new_n399));
  INV_X1    g213(.A(new_n360), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n361), .A2(KEYINPUT81), .A3(G101), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT81), .B1(new_n361), .B2(G101), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n373), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n334), .B(new_n376), .C1(new_n405), .C2(new_n359), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n381), .B2(new_n378), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n399), .B(new_n310), .C1(new_n407), .C2(new_n333), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n398), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT91), .B(new_n311), .C1(new_n384), .C2(new_n397), .ZN(new_n411));
  OAI21_X1  g225(.A(G214), .B1(G237), .B2(G902), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n309), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n288), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(G469), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n323), .B(new_n419), .C1(new_n319), .C2(G128), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT82), .B1(new_n322), .B2(new_n324), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n321), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n340), .A2(new_n343), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n428));
  INV_X1    g242(.A(G134), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(G137), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(G137), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .A3(G134), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n190), .A2(new_n430), .A3(new_n431), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n328), .B1(new_n319), .B2(new_n329), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(new_n372), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n403), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n316), .A2(new_n317), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT67), .B1(new_n319), .B2(new_n313), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n325), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT10), .A3(new_n424), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n427), .A2(new_n438), .A3(new_n441), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT80), .ZN(new_n448));
  INV_X1    g262(.A(G227), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G953), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n448), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n323), .B1(new_n319), .B2(G128), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n318), .B2(new_n320), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n423), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n438), .B1(new_n425), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n457), .B2(KEYINPUT12), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(KEYINPUT12), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n453), .A3(KEYINPUT12), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(KEYINPUT82), .A2(new_n454), .B1(new_n318), .B2(new_n320), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n423), .B1(new_n463), .B2(new_n420), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n441), .B(new_n445), .C1(new_n464), .C2(KEYINPUT10), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n437), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n451), .B1(new_n466), .B2(new_n446), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n292), .B(new_n418), .C1(new_n462), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n425), .A2(new_n456), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT12), .A3(new_n437), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n437), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n461), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n452), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n467), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT86), .A3(new_n418), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n470), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n466), .B1(new_n452), .B2(KEYINPUT84), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n451), .B1(new_n477), .B2(new_n446), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G469), .B1(new_n488), .B2(G902), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n416), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n431), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n429), .A2(G137), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n436), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n436), .A2(KEYINPUT66), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n444), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n439), .A2(KEYINPUT64), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n328), .B(new_n500), .C1(new_n319), .C2(new_n329), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n437), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n444), .A2(new_n436), .A3(new_n493), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n437), .A2(new_n439), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT30), .A4(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(KEYINPUT30), .C1(new_n494), .C2(new_n455), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT68), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n505), .A2(new_n370), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n199), .A2(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n455), .A2(new_n494), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n437), .A2(new_n439), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n370), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT31), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n503), .A2(new_n370), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(KEYINPUT28), .A3(new_n522), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n518), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n512), .A2(new_n533), .A3(new_n518), .A4(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G472), .A2(G902), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT72), .B1(new_n521), .B2(new_n522), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(new_n370), .C1(new_n519), .C2(new_n520), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n523), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT28), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n545), .A2(KEYINPUT29), .A3(new_n518), .A4(new_n527), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n292), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n530), .A2(new_n518), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n512), .A3(new_n523), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT29), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G472), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n539), .A2(new_n540), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n197), .A2(G221), .A3(G234), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT22), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n554), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n560));
  OR3_X1    g374(.A1(new_n559), .A2(new_n432), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n432), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n219), .B1(new_n229), .B2(new_n232), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT74), .B1(new_n312), .B2(G119), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n353), .A3(G128), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n565), .B(new_n567), .C1(new_n353), .C2(G128), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT24), .B(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(KEYINPUT76), .A3(new_n569), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n353), .B2(G128), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n312), .A2(KEYINPUT23), .A3(G119), .ZN(new_n577));
  INV_X1    g391(.A(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n353), .A2(G128), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT75), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n564), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n579), .A3(new_n577), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G110), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n569), .B2(new_n568), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n221), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n563), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(new_n572), .A3(new_n573), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n229), .A2(new_n232), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n219), .A3(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n220), .B(new_n585), .C1(new_n569), .C2(new_n568), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n561), .A4(new_n562), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n593), .A3(new_n292), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT25), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n588), .A2(new_n593), .A3(new_n596), .A4(new_n292), .ZN(new_n597));
  INV_X1    g411(.A(G234), .ZN(new_n598));
  OAI21_X1  g412(.A(G217), .B1(new_n598), .B2(G902), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT73), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n595), .A2(KEYINPUT79), .A3(new_n597), .A4(new_n601), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n601), .A2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n588), .A2(new_n593), .A3(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n414), .A2(new_n490), .A3(new_n552), .A4(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT97), .B(G101), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G3));
  INV_X1    g425(.A(new_n490), .ZN(new_n612));
  INV_X1    g426(.A(new_n537), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n535), .B2(new_n292), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n608), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT98), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n490), .A2(new_n619), .A3(new_n616), .A4(new_n608), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n264), .B1(new_n256), .B2(new_n257), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n287), .A2(new_n290), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n291), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n294), .A2(G902), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n627), .A2(new_n628), .B1(new_n294), .B2(new_n293), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n622), .A2(new_n307), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n398), .A2(new_n408), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n412), .ZN(new_n633));
  INV_X1    g447(.A(new_n412), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT99), .B(new_n634), .C1(new_n398), .C2(new_n408), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n621), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n226), .ZN(G6));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n247), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n188), .B1(new_n237), .B2(new_n246), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT20), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n253), .A2(KEYINPUT102), .A3(new_n187), .A4(new_n188), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n648));
  OR3_X1    g462(.A1(new_n262), .A2(new_n648), .A3(new_n263), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n648), .B1(new_n262), .B2(new_n263), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n298), .A2(new_n647), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n636), .A2(new_n651), .A3(new_n306), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n621), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n591), .A2(new_n592), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n606), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n604), .A2(new_n605), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n662), .A2(new_n613), .A3(new_n615), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n414), .A3(new_n490), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  OR2_X1    g480(.A1(new_n304), .A2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n302), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n490), .A2(new_n651), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n636), .A2(new_n552), .A3(new_n661), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT104), .B(G128), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G30));
  XOR2_X1   g488(.A(new_n668), .B(KEYINPUT39), .Z(new_n675));
  NOR2_X1   g489(.A1(new_n612), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  AOI21_X1  g491(.A(new_n531), .B1(new_n523), .B2(new_n512), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n292), .B1(new_n544), .B2(new_n518), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n539), .A2(new_n540), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n410), .A2(new_n411), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT38), .Z(new_n686));
  INV_X1    g500(.A(new_n298), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n622), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n686), .A2(new_n412), .A3(new_n662), .A4(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n677), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n207), .ZN(G45));
  NOR2_X1   g505(.A1(new_n622), .A2(new_n629), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n490), .A2(new_n692), .A3(new_n668), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n670), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(G146), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G48));
  OAI21_X1  g510(.A(new_n292), .B1(new_n462), .B2(new_n467), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n416), .B1(new_n697), .B2(G469), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT86), .B1(new_n481), .B2(new_n418), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n466), .A2(new_n446), .ZN(new_n700));
  INV_X1    g514(.A(new_n451), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n477), .A2(new_n478), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n702), .A2(new_n469), .A3(G902), .A4(new_n417), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n698), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n698), .B(new_n706), .C1(new_n699), .C2(new_n703), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n705), .A2(KEYINPUT108), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n630), .A2(new_n552), .A3(new_n608), .A4(new_n636), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT41), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G113), .ZN(G15));
  NAND2_X1  g527(.A1(new_n552), .A2(new_n608), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n652), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  INV_X1    g530(.A(new_n707), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n706), .B1(new_n483), .B2(new_n698), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n705), .A2(KEYINPUT108), .A3(new_n707), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n715), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n715), .A2(new_n719), .A3(KEYINPUT109), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  INV_X1    g540(.A(new_n309), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n636), .A3(new_n552), .A4(new_n661), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n705), .A2(new_n707), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n353), .ZN(G21));
  AND2_X1   g545(.A1(new_n545), .A2(new_n527), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n525), .B(new_n534), .C1(new_n732), .C2(new_n518), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n536), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(KEYINPUT110), .A3(new_n536), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n615), .B(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n738), .A2(new_n608), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n688), .A2(new_n636), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n307), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n719), .A3(new_n720), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NAND3_X1  g559(.A1(new_n738), .A2(new_n692), .A3(new_n740), .ZN(new_n746));
  INV_X1    g560(.A(new_n668), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n662), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n705), .A2(new_n748), .A3(new_n636), .A4(new_n707), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n212), .ZN(G27));
  NAND2_X1  g565(.A1(new_n490), .A2(new_n668), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n685), .A2(new_n412), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n552), .A3(new_n608), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n753), .A2(new_n757), .A3(new_n758), .A4(new_n692), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n693), .B2(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(G131), .Z(G33));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n669), .A2(new_n763), .A3(new_n757), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n490), .A2(new_n651), .A3(new_n668), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT112), .B1(new_n765), .B2(new_n756), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n258), .A2(new_n265), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n769), .A2(KEYINPUT43), .A3(new_n629), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT43), .B1(new_n769), .B2(new_n629), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n616), .A2(new_n662), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT44), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n754), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n488), .A2(KEYINPUT45), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n486), .B2(new_n487), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(G469), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n483), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n415), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n675), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n773), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n775), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n791), .A3(new_n415), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n785), .B2(new_n415), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n692), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n608), .A2(new_n747), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n552), .A4(new_n754), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n729), .A2(new_n686), .A3(new_n412), .ZN(new_n802));
  INV_X1    g616(.A(new_n302), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n770), .A2(new_n803), .A3(new_n771), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n804), .A3(new_n741), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT50), .A4(new_n741), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n705), .A2(new_n707), .A3(new_n755), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n608), .A2(new_n803), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n683), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n629), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n769), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n807), .A2(new_n808), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n809), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n804), .A2(KEYINPUT118), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n770), .A2(new_n803), .A3(new_n771), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n809), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n738), .A2(new_n661), .A3(new_n740), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT119), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n824), .B(new_n821), .C1(new_n816), .C2(new_n819), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n814), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n814), .B(KEYINPUT120), .C1(new_n823), .C2(new_n825), .ZN(new_n829));
  INV_X1    g643(.A(G469), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n483), .B1(new_n830), .B2(new_n481), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(new_n415), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n793), .B2(new_n794), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n804), .A2(new_n741), .A3(new_n755), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n814), .B(new_n837), .C1(new_n823), .C2(new_n825), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT116), .B1(new_n793), .B2(new_n794), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n792), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n843), .A3(new_n832), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n839), .B1(new_n844), .B2(new_n834), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n839), .A3(new_n834), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n836), .A2(KEYINPUT51), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n717), .A2(new_n718), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n804), .A2(new_n636), .A3(new_n849), .A4(new_n741), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(new_n300), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n811), .A2(new_n692), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n714), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT48), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n820), .B(new_n856), .C1(KEYINPUT122), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT122), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n801), .B1(new_n848), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n861), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n846), .A2(new_n847), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n826), .A2(new_n827), .B1(new_n834), .B2(new_n833), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n837), .B1(new_n865), .B2(new_n829), .ZN(new_n866));
  OAI211_X1 g680(.A(KEYINPUT123), .B(new_n863), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n609), .B(new_n664), .C1(new_n729), .C2(new_n728), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n711), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n413), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n769), .A3(new_n306), .A4(new_n812), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n769), .A2(new_n687), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n870), .A3(new_n306), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n630), .A2(KEYINPUT113), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n620), .A3(new_n618), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n725), .A2(new_n744), .A3(new_n869), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n490), .A2(new_n748), .A3(new_n755), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n649), .A2(new_n650), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n552), .A2(new_n687), .A3(new_n647), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n746), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n767), .A3(new_n760), .A4(new_n759), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT114), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n711), .ZN(new_n887));
  INV_X1    g701(.A(new_n868), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n878), .A4(new_n744), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n763), .B1(new_n669), .B2(new_n757), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n765), .A2(new_n756), .A3(KEYINPUT112), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n761), .A3(new_n883), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n889), .A2(new_n893), .A3(new_n894), .A4(new_n725), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n746), .A2(new_n749), .ZN(new_n896));
  INV_X1    g710(.A(new_n742), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n683), .A2(new_n753), .A3(new_n662), .A4(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n753), .B(new_n671), .C1(new_n692), .C2(new_n651), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n670), .B1(new_n765), .B2(new_n693), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n750), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT52), .A3(new_n898), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n886), .A2(new_n895), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT53), .ZN(new_n908));
  AND4_X1   g722(.A1(KEYINPUT52), .A2(new_n896), .A3(new_n898), .A4(new_n899), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT52), .B1(new_n904), .B2(new_n898), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT115), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n905), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n895), .A4(new_n886), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n908), .A2(KEYINPUT54), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n907), .A2(new_n915), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n879), .A2(new_n915), .A3(new_n885), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n862), .A2(new_n867), .A3(new_n917), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n299), .A2(new_n197), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n608), .A2(new_n415), .A3(new_n412), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n686), .A2(new_n769), .A3(new_n629), .A4(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n831), .B(KEYINPUT49), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n928), .A3(new_n684), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(G75));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n918), .A2(new_n921), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G902), .ZN(new_n933));
  INV_X1    g747(.A(G210), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n407), .B(new_n333), .Z(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  AND2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n197), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  AOI221_X4 g755(.A(KEYINPUT54), .B1(new_n914), .B2(new_n920), .C1(new_n907), .C2(new_n915), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n919), .B1(new_n918), .B2(new_n921), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n780), .B(KEYINPUT124), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT57), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n944), .A2(new_n946), .B1(new_n462), .B2(new_n467), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n933), .A2(new_n779), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(G54));
  INV_X1    g763(.A(new_n933), .ZN(new_n950));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(new_n253), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n253), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n940), .ZN(G60));
  NAND2_X1  g768(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n922), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n627), .B(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n940), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n917), .A2(new_n922), .ZN(new_n963));
  INV_X1    g777(.A(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n958), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT126), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n942), .B2(new_n943), .ZN(new_n969));
  INV_X1    g783(.A(new_n940), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n588), .A2(new_n593), .ZN(new_n976));
  INV_X1    g790(.A(new_n932), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  INV_X1    g795(.A(new_n659), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n977), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n970), .A4(new_n980), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G66));
  INV_X1    g801(.A(new_n879), .ZN(new_n988));
  AND2_X1   g802(.A1(G224), .A2(G953), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n988), .A2(new_n197), .B1(new_n303), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n407), .B1(G898), .B2(new_n197), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G69));
  NAND3_X1  g806(.A1(new_n505), .A2(new_n509), .A3(new_n511), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(new_n242), .ZN(new_n994));
  INV_X1    g808(.A(new_n690), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n904), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n789), .A2(new_n799), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n996), .B2(KEYINPUT62), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n676), .B(new_n757), .C1(new_n692), .C2(new_n874), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n994), .B1(new_n1001), .B2(new_n197), .ZN(new_n1002));
  INV_X1    g816(.A(G900), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n1003), .B2(new_n197), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n787), .A2(new_n856), .A3(new_n897), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n904), .ZN(new_n1006));
  NOR4_X1   g820(.A1(new_n998), .A2(new_n1006), .A3(new_n761), .A4(new_n892), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1007), .B2(new_n197), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(G953), .B1(new_n449), .B2(new_n1003), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G72));
  INV_X1    g825(.A(new_n678), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  AND3_X1   g828(.A1(new_n1012), .A2(new_n549), .A3(new_n1014), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n908), .A2(new_n916), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1014), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n1007), .B2(new_n988), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n970), .B1(new_n1018), .B2(new_n549), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1014), .B1(new_n1001), .B2(new_n879), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1012), .B1(new_n1020), .B2(KEYINPUT127), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1016), .B(new_n1019), .C1(new_n1021), .C2(new_n1022), .ZN(G57));
endmodule


