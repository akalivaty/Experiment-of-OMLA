//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT92), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT93), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI221_X1 g013(.A(new_n214), .B1(KEYINPUT15), .B2(new_n202), .C1(new_n207), .C2(new_n208), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n207), .A2(new_n213), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n210), .A2(new_n215), .B1(new_n216), .B2(new_n203), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G15gat), .B(G22gat), .Z(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(G1gat), .B1(KEYINPUT95), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n222), .A2(KEYINPUT95), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n226), .B(new_n227), .Z(new_n228));
  NOR2_X1   g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n217), .B(KEYINPUT94), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n218), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n229), .A2(new_n231), .B1(new_n230), .B2(new_n228), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OR3_X1    g033(.A1(new_n234), .A2(KEYINPUT96), .A3(KEYINPUT18), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(new_n228), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n233), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(KEYINPUT96), .B2(KEYINPUT18), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G197gat), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT11), .B(G169gat), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT12), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n247), .A3(new_n239), .A4(new_n238), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G120gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n258), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n257), .A2(new_n259), .A3(G127gat), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT71), .B(G134gat), .C1(new_n258), .C2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n269));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(G169gat), .B2(G176gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n278), .A2(new_n279), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n273), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n282), .A2(new_n279), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(new_n278), .A3(KEYINPUT66), .A4(new_n284), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT25), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  NAND4_X1  g090(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n279), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n294), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(KEYINPUT68), .A3(new_n299), .A4(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n272), .A4(new_n270), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n290), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n281), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n281), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n268), .A2(KEYINPUT26), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n270), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n315), .B(new_n274), .C1(new_n317), .C2(new_n268), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT70), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321));
  AOI211_X1 g120(.A(new_n321), .B(new_n318), .C1(new_n312), .C2(new_n313), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n267), .B1(new_n308), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n282), .B(new_n279), .C1(new_n283), .C2(KEYINPUT65), .ZN(new_n325));
  INV_X1    g124(.A(new_n284), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n286), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n273), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n289), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT69), .B1(new_n301), .B2(new_n303), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n305), .B(new_n302), .C1(new_n296), .C2(new_n300), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n320), .A2(new_n322), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n266), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n337), .B(KEYINPUT64), .Z(new_n338));
  XOR2_X1   g137(.A(G71gat), .B(G99gat), .Z(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n336), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT73), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n336), .A3(new_n338), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(KEYINPUT32), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n324), .A2(new_n336), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n337), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT34), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT34), .ZN(new_n352));
  INV_X1    g151(.A(new_n338), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n345), .B2(new_n347), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n351), .A3(new_n354), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n355), .A4(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT36), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n370));
  XNOR2_X1  g169(.A(G197gat), .B(G204gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT22), .ZN(new_n372));
  INV_X1    g171(.A(G211gat), .ZN(new_n373));
  INV_X1    g172(.A(G218gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G141gat), .B(G148gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(G155gat), .B2(G162gat), .ZN(new_n383));
  OAI221_X1 g182(.A(new_n381), .B1(G155gat), .B2(G162gat), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n381), .B1(G155gat), .B2(G162gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n379), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n387), .A3(new_n370), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n384), .A2(new_n387), .A3(new_n392), .A4(new_n370), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n378), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n401), .B2(new_n388), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n378), .B(KEYINPUT75), .Z(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n399), .B1(new_n398), .B2(new_n404), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  INV_X1    g207(.A(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n398), .A2(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G22gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n414), .B2(new_n405), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n369), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n406), .B2(new_n407), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n412), .A3(new_n405), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n368), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n384), .A2(new_n387), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n260), .B2(new_n265), .ZN(new_n424));
  OAI21_X1  g223(.A(G127gat), .B1(new_n257), .B2(new_n259), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n262), .A2(new_n264), .A3(new_n261), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n388), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n422), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT5), .B1(new_n428), .B2(KEYINPUT82), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n430), .B(new_n422), .C1(new_n424), .C2(new_n427), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT83), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  INV_X1    g232(.A(new_n422), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n425), .A2(new_n388), .A3(new_n426), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n388), .B1(new_n425), .B2(new_n426), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n433), .B1(new_n437), .B2(new_n430), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n428), .A2(KEYINPUT82), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n266), .B1(new_n400), .B2(new_n423), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n391), .A2(new_n393), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n422), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n436), .B(KEYINPUT4), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT0), .ZN(new_n451));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  OAI211_X1 g252(.A(new_n433), .B(new_n422), .C1(new_n443), .C2(new_n444), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n424), .B(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n449), .A2(new_n453), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  INV_X1    g261(.A(new_n453), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n432), .B2(new_n441), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n459), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n453), .B1(new_n449), .B2(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  XOR2_X1   g271(.A(new_n472), .B(KEYINPUT77), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT76), .B1(new_n308), .B2(new_n323), .ZN(new_n475));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(KEYINPUT29), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n334), .A2(new_n479), .A3(new_n335), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n403), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n314), .A2(new_n319), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n334), .A2(new_n483), .A3(new_n477), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n334), .A2(new_n479), .A3(new_n335), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n334), .B2(new_n335), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n477), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n334), .A2(new_n483), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n478), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n378), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n474), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT78), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n476), .B1(new_n475), .B2(new_n480), .ZN(new_n494));
  INV_X1    g293(.A(new_n490), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n395), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n474), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n472), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT30), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n496), .A2(new_n504), .A3(new_n472), .A4(new_n497), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n469), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n502), .A2(KEYINPUT30), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n499), .B1(new_n498), .B2(new_n474), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT78), .B(new_n473), .C1(new_n496), .C2(new_n497), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(KEYINPUT86), .A3(new_n506), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n453), .B(KEYINPUT87), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n456), .A2(new_n458), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n443), .A2(new_n444), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n422), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT39), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n435), .A2(new_n436), .A3(new_n434), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n524), .B2(KEYINPUT88), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(KEYINPUT88), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n529), .A2(KEYINPUT40), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n518), .B1(new_n464), .B2(new_n459), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n529), .B2(KEYINPUT40), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n516), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n459), .B1(new_n442), .B2(new_n448), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT6), .B1(new_n534), .B2(new_n453), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n535), .A2(new_n531), .B1(new_n467), .B2(KEYINPUT6), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n494), .A2(new_n395), .A3(new_n495), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n482), .B1(new_n481), .B2(new_n484), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT37), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT38), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n496), .A2(new_n497), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n474), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n536), .A2(new_n502), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n472), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(KEYINPUT37), .B2(new_n498), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n421), .ZN(new_n551));
  OAI221_X1 g350(.A(new_n367), .B1(new_n421), .B2(new_n507), .C1(new_n533), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT35), .ZN(new_n553));
  AND4_X1   g352(.A1(new_n358), .A2(new_n360), .A3(new_n416), .A4(new_n419), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n507), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n416), .A2(new_n553), .A3(new_n419), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n536), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n501), .A2(KEYINPUT86), .A3(new_n506), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT86), .B1(new_n501), .B2(new_n506), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n364), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n364), .A4(new_n557), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n555), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n250), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G134gat), .ZN(new_n568));
  INV_X1    g367(.A(G162gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT102), .B(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n571), .A2(new_n572), .B1(KEYINPUT8), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT100), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT7), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n575), .B2(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n574), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n231), .A2(new_n219), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n230), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(KEYINPUT103), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(KEYINPUT103), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT104), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n570), .B1(new_n596), .B2(KEYINPUT105), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n592), .A2(new_n594), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n595), .A4(new_n570), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT97), .ZN(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(G57gat), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT98), .A3(G64gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n608), .B(new_n610), .C1(new_n609), .C2(G64gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n614));
  INV_X1    g413(.A(new_n605), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n609), .A2(G64gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n607), .A2(G57gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n604), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n261), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n228), .B1(new_n619), .B2(KEYINPUT21), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G155gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n584), .B(new_n619), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n635), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT106), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n635), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n638), .B2(new_n639), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR4_X1    g449(.A1(new_n636), .A2(new_n642), .A3(new_n646), .A4(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n646), .B1(new_n648), .B2(new_n636), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n633), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n566), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n469), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n224), .ZN(G1324gat));
  INV_X1    g456(.A(new_n516), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n566), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(new_n633), .A3(new_n653), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT16), .B(G8gat), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n222), .B2(new_n660), .ZN(new_n663));
  MUX2_X1   g462(.A(new_n662), .B(new_n663), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g463(.A(G15gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n364), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n655), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT107), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n655), .A2(new_n665), .A3(new_n367), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n421), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n562), .A2(new_n563), .ZN(new_n675));
  INV_X1    g474(.A(new_n555), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(KEYINPUT108), .B(new_n555), .C1(new_n562), .C2(new_n563), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n552), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT109), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n552), .B(new_n681), .C1(new_n677), .C2(new_n678), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n602), .A2(KEYINPUT44), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(KEYINPUT110), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n680), .A2(new_n686), .A3(new_n682), .A4(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n552), .A2(new_n565), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n600), .A2(new_n601), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n469), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n632), .A2(new_n653), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n250), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT111), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n693), .A2(new_n700), .A3(new_n694), .A4(new_n697), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n688), .A2(new_n689), .A3(new_n697), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n469), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT45), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1328gat));
  NOR2_X1   g505(.A1(new_n696), .A2(new_n602), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(G36gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n659), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT112), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(KEYINPUT113), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n685), .A2(new_n692), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n716), .A2(new_n516), .A3(new_n250), .A4(new_n696), .ZN(new_n717));
  OAI221_X1 g516(.A(new_n714), .B1(new_n712), .B2(new_n715), .C1(new_n717), .C2(new_n212), .ZN(G1329gat));
  INV_X1    g517(.A(new_n367), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n719), .B(new_n697), .C1(new_n685), .C2(new_n692), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n708), .A2(G43gat), .A3(new_n666), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n566), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT47), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n723), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n720), .B2(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(KEYINPUT114), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n726), .A2(new_n730), .ZN(G1330gat));
  NOR3_X1   g530(.A1(new_n703), .A2(G50gat), .A3(new_n421), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n420), .B(new_n697), .C1(new_n685), .C2(new_n692), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(G50gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n740), .ZN(G1331gat));
  AND2_X1   g540(.A1(new_n680), .A2(new_n682), .ZN(new_n742));
  INV_X1    g541(.A(new_n653), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n633), .A2(new_n249), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n469), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n609), .ZN(G1332gat));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n658), .A3(new_n744), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n745), .B2(new_n367), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n666), .A2(G71gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n745), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g554(.A1(new_n745), .A2(new_n421), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT116), .B(G78gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n602), .A2(new_n249), .A3(new_n632), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT51), .B1(new_n679), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n759), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n743), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n694), .A3(new_n571), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n249), .A2(new_n743), .A3(new_n632), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n716), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n469), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(new_n571), .ZN(G1336gat));
  AOI21_X1  g569(.A(new_n572), .B1(new_n767), .B2(new_n658), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n516), .A2(G92gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n693), .A2(new_n658), .A3(new_n765), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n768), .B2(new_n367), .ZN(new_n781));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n782), .A3(new_n364), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1338gat));
  XNOR2_X1  g583(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n767), .B2(new_n420), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n421), .A2(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n763), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n693), .A2(new_n420), .A3(new_n765), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n790), .A3(new_n785), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(new_n632), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n232), .A2(new_n233), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n236), .A2(new_n237), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n244), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n248), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT54), .B1(new_n640), .B2(new_n635), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n642), .A2(new_n650), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n646), .B1(new_n641), .B2(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n642), .A2(new_n802), .A3(new_n650), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n804), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n651), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n806), .A2(new_n809), .A3(new_n651), .A4(KEYINPUT118), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n689), .A2(new_n801), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n249), .A3(new_n813), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n801), .A2(new_n653), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n689), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n797), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n654), .A2(new_n250), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT119), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n469), .A3(new_n658), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n554), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(KEYINPUT120), .A3(new_n554), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n253), .A3(new_n249), .ZN(new_n831));
  INV_X1    g630(.A(new_n823), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n822), .B1(new_n818), .B2(new_n819), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n658), .A2(new_n469), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n666), .A2(new_n420), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n250), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n838), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n251), .A3(new_n653), .ZN(new_n840));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837), .B2(new_n743), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1341gat));
  XOR2_X1   g641(.A(KEYINPUT71), .B(G127gat), .Z(new_n843));
  NOR3_X1   g642(.A1(new_n837), .A2(new_n797), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n554), .A3(new_n632), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n843), .ZN(G1342gat));
  NOR2_X1   g645(.A1(new_n602), .A2(G134gat), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n826), .A2(KEYINPUT56), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n837), .B2(new_n602), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT56), .B1(new_n826), .B2(new_n848), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n719), .A2(new_n421), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n821), .A2(new_n694), .A3(new_n823), .A4(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT121), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n250), .A2(G141gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT121), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n855), .A2(new_n516), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n821), .A2(new_n420), .A3(new_n823), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n250), .A2(new_n810), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n689), .B1(new_n862), .B2(new_n816), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n797), .B1(new_n863), .B2(new_n814), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n819), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n421), .A2(new_n861), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n860), .A2(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n835), .A2(new_n367), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n250), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(G141gat), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n858), .B(new_n859), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n825), .A2(new_n853), .A3(new_n856), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n867), .A2(new_n250), .A3(new_n868), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n867), .A2(new_n868), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n877), .C1(new_n878), .C2(new_n653), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n880));
  AND3_X1   g679(.A1(new_n821), .A2(new_n823), .A3(new_n866), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n689), .A2(new_n801), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n810), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n797), .B1(new_n863), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n819), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n885), .B2(new_n420), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n868), .A2(new_n743), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n880), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n855), .A2(new_n516), .A3(new_n857), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n653), .A2(new_n877), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n879), .A2(new_n890), .B1(new_n891), .B2(new_n892), .ZN(G1345gat));
  NOR3_X1   g692(.A1(new_n867), .A2(new_n797), .A3(new_n868), .ZN(new_n894));
  INV_X1    g693(.A(G155gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n632), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n894), .A2(new_n895), .B1(new_n891), .B2(new_n896), .ZN(G1346gat));
  OR2_X1    g696(.A1(new_n891), .A2(new_n602), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n602), .A2(new_n569), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n898), .A2(new_n569), .B1(new_n878), .B2(new_n899), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n516), .A2(new_n694), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n834), .A2(new_n836), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n250), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n834), .A2(new_n554), .A3(new_n901), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n249), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(G1348gat));
  INV_X1    g708(.A(G176gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n653), .ZN(new_n911));
  OAI21_X1  g710(.A(G176gat), .B1(new_n902), .B2(new_n743), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n309), .A3(new_n632), .ZN(new_n914));
  OAI21_X1  g713(.A(G183gat), .B1(new_n902), .B2(new_n797), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n904), .A2(new_n281), .A3(new_n689), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n902), .B2(new_n602), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(G190gat), .C1(new_n902), .C2(new_n602), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n918), .B1(new_n920), .B2(new_n923), .ZN(G1351gat));
  AND2_X1   g723(.A1(new_n367), .A2(new_n901), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n834), .A2(new_n420), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n250), .A2(G197gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT125), .Z(new_n929));
  NAND2_X1  g728(.A1(new_n887), .A2(new_n925), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n250), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1352gat));
  OAI21_X1  g731(.A(G204gat), .B1(new_n930), .B2(new_n743), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n743), .A2(G204gat), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n926), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n933), .B(new_n935), .C1(new_n938), .C2(new_n939), .ZN(G1353gat));
  OAI211_X1 g739(.A(new_n632), .B(new_n925), .C1(new_n881), .C2(new_n886), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n632), .A2(new_n373), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n942), .A2(new_n943), .B1(new_n926), .B2(new_n944), .ZN(G1354gat));
  OAI21_X1  g744(.A(G218gat), .B1(new_n930), .B2(new_n602), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n689), .A2(new_n374), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n926), .B2(new_n947), .ZN(G1355gat));
endmodule


