//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G107), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT82), .A3(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n193), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(G104), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n191), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G101), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT83), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT83), .A2(G101), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n191), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n204), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT2), .B(G113), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G116), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n214), .A2(new_n216), .A3(G119), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT67), .B1(new_n213), .B2(G119), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n212), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT2), .B(G113), .Z(new_n224));
  NAND3_X1  g038(.A1(new_n214), .A2(new_n216), .A3(G119), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n218), .A4(new_n221), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(KEYINPUT69), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(new_n212), .C1(new_n217), .C2(new_n222), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n189), .B1(new_n211), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G110), .B(G122), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n207), .B1(new_n196), .B2(new_n197), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n233), .A2(new_n199), .B1(new_n198), .B2(new_n200), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n203), .A2(KEYINPUT4), .A3(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n236), .A2(KEYINPUT88), .A3(new_n229), .A4(new_n227), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT84), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n190), .B2(G107), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n193), .A2(KEYINPUT84), .A3(G104), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n191), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G101), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT86), .B1(new_n243), .B2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n209), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n217), .A2(new_n222), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n213), .A2(KEYINPUT5), .A3(G119), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n249), .A2(new_n252), .B1(new_n224), .B2(new_n248), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n231), .A2(new_n232), .A3(new_n237), .A4(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n231), .A2(new_n254), .A3(new_n237), .ZN(new_n258));
  INV_X1    g072(.A(new_n232), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  INV_X1    g081(.A(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G143), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n269), .B2(KEYINPUT1), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n265), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n266), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n269), .A2(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n269), .A2(new_n271), .A3(new_n278), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n264), .B(new_n275), .C1(new_n281), .C2(new_n265), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n279), .A2(new_n280), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT90), .A3(G125), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G224), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G953), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n285), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n263), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n247), .A2(new_n253), .A3(KEYINPUT91), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n232), .B(KEYINPUT8), .ZN(new_n293));
  INV_X1    g107(.A(new_n254), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n202), .A2(new_n208), .B1(G101), .B2(new_n241), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n253), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n285), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n300), .B2(new_n287), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n285), .A2(new_n299), .A3(KEYINPUT7), .A4(new_n288), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n304), .B2(new_n255), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n290), .A2(new_n291), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n291), .ZN(new_n307));
  INV_X1    g121(.A(new_n289), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n261), .B2(new_n262), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n311));
  INV_X1    g125(.A(new_n255), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n188), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  OAI21_X1  g130(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT81), .Z(new_n318));
  INV_X1    g132(.A(G469), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT73), .B(G902), .Z(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(G227), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT1), .B1(new_n270), .B2(G146), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n327), .A2(G128), .B1(new_n269), .B2(new_n271), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT70), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(KEYINPUT10), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n244), .B2(new_n246), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n334));
  OAI21_X1  g148(.A(G128), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(G143), .B2(new_n268), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT85), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n272), .B1(new_n339), .B2(new_n274), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT10), .B1(new_n340), .B2(new_n296), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n283), .B1(new_n234), .B2(new_n235), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n333), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G134), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT11), .B1(new_n344), .B2(G137), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT11), .ZN(new_n346));
  INV_X1    g160(.A(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT65), .B1(new_n347), .B2(G134), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT65), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n344), .A3(G137), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT64), .A2(G131), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT64), .A2(G131), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n349), .A2(new_n350), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n350), .A2(new_n352), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n349), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT87), .B1(new_n343), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n332), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n247), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n236), .A2(new_n281), .ZN(new_n365));
  INV_X1    g179(.A(new_n335), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n327), .A2(new_n334), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n274), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n296), .B1(new_n368), .B2(new_n329), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n364), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n373));
  INV_X1    g187(.A(new_n361), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n362), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n364), .A2(new_n365), .A3(new_n371), .A4(new_n361), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n325), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n244), .A2(new_n380), .A3(new_n246), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n369), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT12), .B1(new_n382), .B2(new_n374), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT12), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n384), .B(new_n361), .C1(new_n381), .C2(new_n369), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n325), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n319), .B(new_n320), .C1(new_n378), .C2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n319), .A2(new_n310), .ZN(new_n390));
  INV_X1    g204(.A(new_n387), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n377), .B1(new_n383), .B2(new_n385), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n376), .A2(new_n391), .B1(new_n392), .B2(new_n324), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n393), .B2(G469), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n318), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(new_n268), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n268), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G237), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n322), .A3(G214), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n270), .ZN(new_n404));
  NOR2_X1   g218(.A1(G237), .A2(G953), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(G143), .A3(G214), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n399), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n406), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT94), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT94), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n415), .B(new_n400), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n190), .ZN(new_n419));
  INV_X1    g233(.A(G140), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G125), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n265), .A2(G140), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT16), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n265), .A2(KEYINPUT16), .A3(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n268), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n424), .A3(G146), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n355), .B1(new_n404), .B2(new_n406), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n404), .A2(new_n355), .A3(new_n406), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n430), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT95), .B1(new_n430), .B2(KEYINPUT17), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n429), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n417), .A2(new_n419), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n419), .B1(new_n417), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n310), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G475), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n419), .ZN(new_n444));
  INV_X1    g258(.A(new_n412), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT93), .B1(new_n404), .B2(new_n406), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n401), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n415), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n413), .A2(KEYINPUT94), .A3(new_n401), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n408), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n427), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n431), .A2(new_n433), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n396), .B(KEYINPUT19), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n268), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT79), .A4(G146), .ZN(new_n456));
  AND4_X1   g270(.A1(new_n452), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n444), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n417), .A2(new_n419), .A3(new_n437), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n443), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND4_X1   g279(.A1(KEYINPUT96), .A2(new_n461), .A3(new_n464), .A4(new_n442), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n441), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G952), .ZN(new_n468));
  AOI211_X1 g282(.A(G953), .B(new_n468), .C1(G234), .C2(G237), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n322), .B(new_n320), .C1(G234), .C2(G237), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G898), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n214), .A2(new_n216), .A3(G122), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n213), .A2(G122), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT14), .A4(G122), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(G107), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n193), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n270), .A2(G128), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n266), .B2(G143), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n270), .A2(KEYINPUT97), .A3(G128), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G134), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT97), .B1(new_n270), .B2(G128), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n266), .A3(G143), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n344), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n478), .B(new_n479), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT13), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n484), .A3(G134), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n488), .B(new_n480), .C1(new_n491), .C2(new_n344), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n193), .B1(new_n473), .B2(new_n475), .ZN(new_n495));
  INV_X1    g309(.A(new_n479), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G217), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n316), .A2(new_n498), .A3(G953), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n490), .B2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n320), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n504), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n467), .A2(new_n472), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n315), .A2(new_n395), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n498), .B1(new_n320), .B2(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT22), .B(G137), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT80), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n220), .A2(G128), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n266), .A2(G119), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT74), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n266), .A2(G119), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n220), .A2(G128), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT75), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n518), .A2(new_n526), .A3(new_n522), .A4(new_n523), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n428), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT76), .B1(new_n266), .B2(G119), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT76), .B(KEYINPUT23), .C1(new_n266), .C2(G119), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT77), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT23), .B1(new_n516), .B2(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n520), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n533), .A2(G110), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n515), .B1(new_n528), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n426), .A2(new_n427), .B1(new_n524), .B2(KEYINPUT75), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n533), .A2(G110), .A3(new_n537), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(KEYINPUT78), .A3(new_n541), .A4(new_n527), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n452), .A2(new_n456), .A3(new_n398), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n531), .A2(G110), .A3(new_n532), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n523), .B1(new_n518), .B2(new_n522), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n514), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n548), .B(new_n513), .C1(new_n539), .C2(new_n542), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT25), .B1(new_n552), .B2(new_n320), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n554));
  INV_X1    g368(.A(new_n320), .ZN(new_n555));
  NOR4_X1   g369(.A1(new_n550), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n510), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n510), .A2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n552), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n281), .B1(new_n357), .B2(new_n360), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT66), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n344), .B2(G137), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n344), .A2(G137), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n347), .A2(KEYINPUT66), .A3(G134), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G131), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n330), .A2(new_n356), .A3(new_n570), .A4(new_n331), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n571), .A3(KEYINPUT30), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n345), .A2(new_n348), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n350), .A2(new_n352), .ZN(new_n575));
  OAI21_X1  g389(.A(G131), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n283), .B1(new_n576), .B2(new_n356), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n356), .A2(new_n379), .A3(new_n570), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n227), .A2(new_n229), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n572), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n230), .A2(new_n564), .A3(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n405), .A2(G210), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT27), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT26), .B(G101), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT31), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n586), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n564), .A2(new_n571), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT28), .B1(new_n590), .B2(new_n230), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n230), .A2(KEYINPUT28), .A3(new_n564), .A4(new_n571), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n229), .B(new_n227), .C1(new_n577), .C2(new_n578), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n589), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n572), .A2(new_n579), .A3(new_n580), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT31), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n586), .A4(new_n582), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n588), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT71), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n588), .A2(new_n595), .A3(new_n598), .A4(KEYINPUT71), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n563), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT32), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n602), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n562), .A2(KEYINPUT32), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT29), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n592), .A2(new_n593), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT28), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n582), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n589), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n596), .A2(new_n589), .A3(new_n582), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n582), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n564), .A2(new_n571), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n580), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n230), .A2(KEYINPUT72), .A3(new_n564), .A4(new_n571), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT28), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(KEYINPUT29), .A3(new_n586), .A4(new_n611), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n614), .A2(new_n622), .A3(new_n320), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n606), .A2(new_n607), .B1(new_n623), .B2(G472), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n561), .B1(new_n605), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n509), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n205), .A2(new_n206), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G3));
  INV_X1    g442(.A(new_n510), .ZN(new_n629));
  INV_X1    g443(.A(new_n513), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n543), .A2(new_n549), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n548), .B1(new_n539), .B2(new_n542), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n631), .B(new_n320), .C1(new_n632), .C2(new_n514), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n554), .ZN(new_n634));
  INV_X1    g448(.A(new_n550), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(KEYINPUT25), .A3(new_n320), .A4(new_n631), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n629), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n558), .B2(new_n552), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n395), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n603), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n555), .B1(new_n601), .B2(new_n602), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n306), .A2(new_n314), .ZN(new_n647));
  INV_X1    g461(.A(new_n472), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n187), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n490), .A2(new_n497), .ZN(new_n650));
  INV_X1    g464(.A(new_n499), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n503), .A3(new_n320), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT33), .B1(new_n500), .B2(new_n501), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n652), .A2(new_n657), .A3(new_n653), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n555), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n655), .B1(new_n659), .B2(new_n503), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT99), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(new_n655), .C1(new_n659), .C2(new_n503), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n467), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n649), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n646), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  XNOR2_X1  g483(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n440), .A2(G475), .B1(new_n460), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n461), .A2(new_n442), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n507), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n315), .A2(new_n648), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n646), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  INV_X1    g494(.A(new_n632), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT36), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n514), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n632), .B1(new_n682), .B2(new_n514), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n684), .A2(new_n685), .A3(new_n559), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT101), .B1(new_n557), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n637), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n643), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n509), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT102), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  INV_X1    g509(.A(G900), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n469), .B1(new_n470), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n672), .A2(new_n507), .A3(new_n674), .A4(new_n698), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n188), .B(new_n699), .C1(new_n306), .C2(new_n314), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n688), .A2(new_n690), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n606), .A2(new_n607), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n623), .A2(G472), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n702), .B(new_n703), .C1(KEYINPUT32), .C2(new_n603), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n395), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  INV_X1    g520(.A(KEYINPUT38), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n647), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n634), .A2(new_n636), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n686), .B1(new_n709), .B2(new_n510), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n507), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT96), .B1(new_n458), .B2(new_n459), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n673), .B1(new_n713), .B2(KEYINPUT20), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n463), .A2(new_n460), .A3(new_n464), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n712), .B1(new_n716), .B2(new_n441), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n310), .B1(new_n620), .B2(new_n586), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n589), .B1(new_n596), .B2(new_n582), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n702), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n717), .B1(new_n721), .B2(new_n604), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n708), .A2(new_n188), .A3(new_n711), .A4(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n697), .B(KEYINPUT39), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n395), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT40), .Z(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  OAI21_X1  g544(.A(new_n689), .B1(new_n637), .B2(new_n686), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n710), .A2(KEYINPUT101), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n704), .A2(new_n395), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n664), .A2(new_n467), .A3(new_n698), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n315), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n268), .ZN(G48));
  AND3_X1   g552(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n377), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n388), .B1(new_n741), .B2(new_n324), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(new_n555), .ZN(new_n743));
  INV_X1    g557(.A(new_n318), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n389), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n666), .A2(new_n625), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n677), .A2(new_n625), .A3(new_n745), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT104), .B(G116), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G18));
  AND4_X1   g565(.A1(new_n704), .A2(new_n508), .A3(new_n731), .A4(new_n732), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n647), .A2(new_n187), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n743), .A2(new_n744), .A3(new_n389), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  NAND4_X1  g571(.A1(new_n717), .A2(new_n743), .A3(new_n744), .A4(new_n389), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n649), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n588), .A2(new_n598), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n621), .A2(new_n611), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n586), .B1(new_n761), .B2(KEYINPUT105), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n621), .A2(new_n763), .A3(new_n611), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  OAI22_X1  g579(.A1(new_n765), .A2(new_n563), .B1(new_n642), .B2(new_n641), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n561), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NOR2_X1   g583(.A1(new_n642), .A2(new_n641), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n618), .A2(new_n619), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n610), .B1(new_n771), .B2(new_n616), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT105), .B1(new_n772), .B2(new_n591), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n589), .A3(new_n764), .ZN(new_n774));
  INV_X1    g588(.A(new_n760), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n563), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n770), .A2(new_n776), .A3(new_n710), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n315), .A3(new_n735), .A4(new_n745), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  NOR2_X1   g593(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n306), .A2(new_n187), .A3(new_n314), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n704), .A3(new_n638), .A4(new_n395), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n782), .B2(new_n734), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n389), .A2(new_n394), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n744), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n306), .A2(new_n187), .A3(new_n314), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n780), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n625), .A3(new_n735), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  INV_X1    g605(.A(new_n699), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n625), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  NAND2_X1  g608(.A1(new_n393), .A2(KEYINPUT45), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n392), .A2(new_n324), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n387), .B1(new_n362), .B2(new_n375), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n799), .A3(G469), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n795), .A2(new_n799), .A3(KEYINPUT107), .A4(G469), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n390), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n389), .B1(new_n804), .B2(KEYINPUT46), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n806), .B(new_n390), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n744), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(new_n726), .ZN(new_n810));
  INV_X1    g624(.A(new_n467), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT43), .B1(new_n811), .B2(KEYINPUT108), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n664), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n811), .B(new_n664), .C1(KEYINPUT108), .C2(KEYINPUT43), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n643), .A3(new_n711), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n819), .A2(new_n820), .A3(new_n786), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT109), .B(G137), .Z(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G39));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n808), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT47), .B(new_n744), .C1(new_n805), .C2(new_n807), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n704), .A2(new_n786), .A3(new_n638), .A4(new_n734), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  AND2_X1   g645(.A1(new_n743), .A2(new_n389), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n318), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n827), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n469), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n814), .B2(new_n815), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(new_n767), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n781), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n754), .A2(new_n786), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n777), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n721), .A2(new_n604), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n638), .A3(new_n469), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n745), .A2(new_n781), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT118), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n561), .A2(new_n835), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n840), .A2(new_n846), .A3(new_n842), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n664), .A2(new_n467), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n841), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n754), .A2(new_n187), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n708), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n767), .A3(new_n836), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n708), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n857), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n837), .A3(KEYINPUT50), .A4(new_n855), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT51), .B1(new_n839), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n468), .B(G953), .C1(new_n837), .C2(new_n755), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n836), .A2(new_n625), .A3(new_n840), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n865));
  XNOR2_X1  g679(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n863), .B(new_n866), .C1(new_n665), .C2(new_n849), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n839), .A2(new_n861), .A3(KEYINPUT51), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n839), .A2(new_n861), .A3(new_n870), .A4(KEYINPUT51), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n862), .B(new_n867), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n873));
  AND4_X1   g687(.A1(new_n704), .A2(new_n395), .A3(new_n731), .A4(new_n732), .ZN(new_n874));
  INV_X1    g688(.A(new_n736), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n637), .A2(new_n686), .A3(new_n697), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n315), .A2(new_n395), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n722), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n874), .A2(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n766), .A2(new_n734), .A3(new_n710), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n874), .A2(new_n700), .B1(new_n755), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT112), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n705), .A2(new_n778), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n315), .A2(new_n395), .A3(new_n876), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n733), .A2(new_n736), .B1(new_n885), .B2(new_n722), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(KEYINPUT52), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n625), .B(new_n745), .C1(new_n666), .C2(new_n677), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n755), .A2(new_n752), .B1(new_n759), .B2(new_n767), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n790), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n665), .A2(KEYINPUT110), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n664), .A2(new_n467), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n892), .B(new_n894), .C1(new_n467), .C2(new_n712), .ZN(new_n895));
  INV_X1    g709(.A(new_n649), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n644), .A4(new_n639), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n509), .B1(new_n691), .B2(new_n625), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n675), .A2(new_n712), .A3(new_n698), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n787), .A2(new_n704), .A3(new_n701), .A4(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n793), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT111), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n770), .A2(new_n776), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n735), .A3(new_n711), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n781), .A2(new_n395), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n787), .A3(KEYINPUT111), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n888), .A2(new_n891), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(new_n882), .B2(new_n887), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n873), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n790), .A2(new_n890), .A3(KEYINPUT53), .A4(new_n889), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n900), .A2(new_n793), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n906), .A2(new_n907), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n897), .A4(new_n898), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n916), .B2(KEYINPUT116), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n882), .A2(new_n887), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT52), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT52), .B1(new_n884), .B2(new_n886), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n917), .A2(new_n920), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n923), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n909), .A2(new_n891), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT113), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT113), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n933), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n910), .A2(new_n873), .A3(new_n911), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n790), .A2(new_n889), .A3(new_n890), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n916), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n920), .A2(new_n939), .A3(new_n888), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT115), .B1(new_n940), .B2(new_n873), .ZN(new_n941));
  AOI22_X1  g755(.A1(new_n932), .A2(new_n934), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n872), .B(new_n927), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n468), .A2(new_n322), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n832), .B(KEYINPUT49), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n813), .A2(new_n561), .A3(new_n318), .A4(new_n188), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n947), .A2(new_n842), .A3(new_n708), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(G75));
  NOR2_X1   g764(.A1(new_n322), .A2(G952), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n320), .B1(new_n912), .B2(new_n924), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT56), .B1(new_n953), .B2(new_n307), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n263), .A2(new_n289), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n309), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT55), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n952), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n320), .B(new_n291), .C1(new_n912), .C2(new_n924), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n960), .A2(KEYINPUT56), .A3(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT121), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n954), .A2(new_n958), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n960), .B2(KEYINPUT56), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n952), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n966), .ZN(G51));
  XNOR2_X1  g781(.A(new_n925), .B(new_n943), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n390), .B(KEYINPUT122), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT57), .ZN(new_n970));
  OAI22_X1  g784(.A1(new_n968), .A2(new_n970), .B1(new_n378), .B2(new_n388), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n953), .A2(new_n802), .A3(new_n803), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n951), .B1(new_n971), .B2(new_n972), .ZN(G54));
  AND3_X1   g787(.A1(new_n953), .A2(KEYINPUT58), .A3(G475), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n952), .B1(new_n974), .B2(new_n461), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n461), .B2(new_n974), .ZN(G60));
  NAND2_X1  g790(.A1(new_n656), .A2(new_n658), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT59), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n952), .B1(new_n968), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n932), .A2(new_n934), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n937), .A2(new_n941), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n943), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n985), .B2(new_n926), .ZN(new_n986));
  INV_X1    g800(.A(new_n977), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(G63));
  NOR2_X1   g802(.A1(new_n684), .A2(new_n685), .ZN(new_n989));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT60), .Z(new_n991));
  NAND3_X1  g805(.A1(new_n925), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n925), .A2(new_n991), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n952), .B(new_n992), .C1(new_n993), .C2(new_n552), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT61), .B1(new_n992), .B2(KEYINPUT123), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G66));
  OAI21_X1  g810(.A(G953), .B1(new_n471), .B2(new_n286), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n890), .A2(new_n889), .A3(new_n897), .A4(new_n898), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n322), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n261), .B(new_n262), .C1(G898), .C2(new_n322), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1000), .B(new_n1001), .Z(G69));
  NOR2_X1   g816(.A1(new_n884), .A2(new_n737), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n729), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1005), .A2(new_n729), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n895), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n625), .A2(new_n781), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n727), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n810), .B2(new_n821), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1007), .A2(new_n830), .A3(new_n1009), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n322), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n572), .A2(new_n579), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(new_n454), .Z(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(G900), .B2(G953), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n810), .A2(new_n625), .A3(new_n315), .A4(new_n717), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(new_n822), .A3(new_n1005), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT126), .B1(new_n790), .B2(new_n793), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n790), .A2(KEYINPUT126), .A3(new_n793), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n830), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1020), .B1(new_n1026), .B2(G953), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1029), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1019), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(G72));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  OAI21_X1  g849(.A(new_n1035), .B1(new_n1014), .B2(new_n999), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n719), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1022), .A2(new_n1025), .A3(new_n999), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1035), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n613), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1037), .A2(new_n1040), .A3(new_n952), .ZN(new_n1041));
  NOR4_X1   g855(.A1(new_n942), .A2(new_n613), .A3(new_n719), .A4(new_n1039), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(G57));
endmodule


