//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT86), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT90), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n214), .B1(new_n213), .B2(new_n215), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n208), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n218), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT92), .A3(new_n216), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT14), .B(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G29gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229));
  INV_X1    g028(.A(G50gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(G43gat), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G43gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G50gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n222), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n233), .A2(KEYINPUT87), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(G43gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT87), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n236), .A2(KEYINPUT88), .A3(new_n238), .A4(new_n229), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n225), .A2(new_n227), .B1(new_n233), .B2(new_n231), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n235), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n225), .A2(new_n227), .ZN(new_n246));
  INV_X1    g045(.A(new_n234), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT89), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n219), .A2(new_n221), .A3(new_n244), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(KEYINPUT17), .A3(new_n244), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n217), .A2(new_n218), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT91), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n249), .A2(KEYINPUT17), .A3(new_n244), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT17), .B1(new_n249), .B2(new_n244), .ZN(new_n262));
  OAI211_X1 g061(.A(KEYINPUT91), .B(new_n259), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT18), .B(new_n253), .C1(new_n260), .C2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n251), .B(KEYINPUT13), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n219), .A2(new_n221), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n254), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n269), .B2(new_n250), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n263), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n278), .B2(new_n253), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n207), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n252), .B1(new_n277), .B2(new_n263), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n270), .B1(new_n281), .B2(KEYINPUT18), .ZN(new_n282));
  INV_X1    g081(.A(new_n206), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n253), .B1(new_n260), .B2(new_n264), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n273), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  INV_X1    g090(.A(G155gat), .ZN(new_n292));
  INV_X1    g091(.A(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(KEYINPUT2), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G141gat), .B(G148gat), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n295), .B(new_n294), .C1(new_n299), .C2(KEYINPUT2), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g102(.A1(G211gat), .A2(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307));
  AND2_X1   g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n303), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT3), .B1(new_n315), .B2(KEYINPUT80), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n310), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n313), .A3(new_n306), .ZN(new_n318));
  AOI211_X1 g117(.A(KEYINPUT80), .B(KEYINPUT29), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n302), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n298), .A2(new_n300), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n314), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G228gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n290), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n317), .B2(new_n318), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n301), .B1(new_n336), .B2(new_n319), .ZN(new_n337));
  INV_X1    g136(.A(new_n331), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n326), .B2(new_n327), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(KEYINPUT81), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n322), .B1(new_n327), .B2(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n301), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n331), .B1(new_n343), .B2(new_n328), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n289), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g145(.A(G22gat), .B(new_n344), .C1(new_n333), .C2(new_n340), .ZN(new_n347));
  OAI21_X1  g146(.A(G78gat), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n340), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT81), .B1(new_n337), .B2(new_n339), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G22gat), .ZN(new_n352));
  INV_X1    g151(.A(G78gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n341), .A2(new_n289), .A3(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT31), .B(G50gat), .ZN(new_n356));
  INV_X1    g155(.A(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n348), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n348), .B2(new_n355), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G15gat), .B(G43gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT74), .ZN(new_n364));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT64), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT24), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(KEYINPUT23), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n371), .A2(new_n376), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n383));
  INV_X1    g182(.A(G176gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n383), .A2(KEYINPUT23), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT67), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G169gat), .A3(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(KEYINPUT28), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399));
  OR2_X1    g198(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n378), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT26), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT68), .B1(G169gat), .B2(G176gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT71), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT71), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n378), .B2(new_n409), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n392), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n372), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n394), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n396), .A3(new_n401), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n376), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT70), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n376), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n379), .A2(new_n381), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n408), .A2(KEYINPUT23), .A3(new_n410), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n392), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n387), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G113gat), .B(G120gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n429), .B2(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n417), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  INV_X1    g239(.A(new_n372), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n392), .A2(new_n412), .A3(new_n414), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(new_n411), .ZN(new_n443));
  AND2_X1   g242(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT27), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n403), .ZN(new_n447));
  AOI21_X1  g246(.A(G190gat), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n397), .B1(new_n448), .B2(KEYINPUT28), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n443), .A2(new_n449), .B1(new_n393), .B2(new_n382), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n418), .A2(new_n376), .A3(new_n421), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n421), .B1(new_n418), .B2(new_n376), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT25), .B1(new_n453), .B2(new_n426), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n440), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n368), .B1(new_n439), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n366), .B1(new_n456), .B2(KEYINPUT32), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(KEYINPUT73), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT73), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n438), .B1(new_n417), .B2(new_n428), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(new_n440), .A3(new_n454), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n367), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(KEYINPUT33), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT75), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n366), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n366), .A2(new_n466), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT33), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n456), .B(KEYINPUT32), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(KEYINPUT77), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n462), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n368), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n479), .A3(new_n477), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n473), .A2(new_n474), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n482), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n485), .A2(new_n480), .B1(new_n477), .B2(new_n476), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(KEYINPUT77), .A3(new_n470), .A4(new_n465), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n362), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n417), .A2(new_n428), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n496), .B2(new_n325), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n493), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n327), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  INV_X1    g299(.A(new_n327), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n495), .A2(KEYINPUT29), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n494), .ZN(new_n503));
  XNOR2_X1  g302(.A(G8gat), .B(G36gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(G64gat), .B(G92gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n499), .A2(new_n503), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT30), .A4(new_n506), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n435), .A2(new_n437), .A3(new_n298), .A4(new_n300), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n435), .A2(new_n437), .B1(new_n298), .B2(new_n300), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n323), .A3(new_n438), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n524), .A3(new_n515), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  XNOR2_X1  g329(.A(G1gat), .B(G29gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT0), .ZN(new_n532));
  XOR2_X1   g331(.A(G57gat), .B(G85gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT6), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n541), .A3(new_n536), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT84), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(KEYINPUT84), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n514), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n492), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n488), .A2(new_n549), .A3(new_n361), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n488), .B2(new_n361), .ZN(new_n551));
  INV_X1    g350(.A(new_n514), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n535), .B1(new_n536), .B2(KEYINPUT79), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n540), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n557), .B2(new_n544), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT38), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n511), .B1(new_n510), .B2(KEYINPUT37), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n510), .A2(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n538), .A2(new_n540), .A3(new_n507), .A4(new_n542), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n500), .B(new_n327), .C1(new_n502), .C2(new_n494), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n501), .B1(new_n497), .B2(new_n498), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT37), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n560), .A2(new_n568), .A3(KEYINPUT38), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n517), .B(KEYINPUT4), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n515), .B1(new_n571), .B2(new_n524), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n518), .A2(new_n519), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT39), .B1(new_n573), .B2(new_n516), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT39), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n534), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT40), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n514), .A2(new_n535), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n361), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n556), .ZN(new_n584));
  OAI22_X1  g383(.A1(new_n570), .A2(new_n583), .B1(new_n584), .B2(new_n361), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n484), .A2(KEYINPUT36), .A3(new_n487), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT36), .B1(new_n484), .B2(new_n487), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n288), .B1(new_n558), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G134gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G162gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G99gat), .B(G106gat), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n601), .A3(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n254), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n593), .A2(new_n594), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n611), .B1(new_n261), .B2(new_n262), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n599), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n597), .B1(new_n616), .B2(KEYINPUT96), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n598), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n615), .A3(new_n599), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT96), .A4(new_n597), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G71gat), .B(G78gat), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n627));
  XOR2_X1   g426(.A(G57gat), .B(G64gat), .Z(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G71gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n353), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(KEYINPUT9), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI221_X1 g432(.A(new_n628), .B1(KEYINPUT9), .B2(new_n631), .C1(new_n626), .C2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT21), .ZN(new_n636));
  XNOR2_X1  g435(.A(G127gat), .B(G155gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n219), .A2(new_n221), .B1(KEYINPUT21), .B2(new_n635), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT95), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n640), .B(new_n646), .Z(new_n647));
  NOR2_X1   g446(.A1(new_n625), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n611), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n635), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n611), .A2(new_n634), .A3(new_n633), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(KEYINPUT97), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n650), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n649), .A2(KEYINPUT10), .A3(new_n635), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(KEYINPUT97), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n656), .A2(new_n661), .A3(new_n666), .A4(new_n662), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n592), .A2(new_n648), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n555), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n211), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n552), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n678), .B(new_n679), .C1(new_n214), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n588), .B2(new_n589), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n488), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT98), .A3(new_n587), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n672), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n490), .A2(new_n491), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n672), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n361), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  INV_X1    g494(.A(new_n474), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT77), .B1(new_n465), .B2(new_n470), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(new_n697), .A3(new_n486), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n483), .A2(new_n471), .A3(new_n472), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n361), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT85), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n488), .A2(new_n549), .A3(new_n361), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n584), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT35), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n704), .A2(new_n548), .B1(new_n586), .B2(new_n686), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n695), .B1(new_n705), .B2(new_n624), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n703), .A2(KEYINPUT35), .B1(new_n492), .B2(new_n547), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n625), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n647), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n670), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n287), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n555), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n625), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT99), .Z(new_n717));
  OAI211_X1 g516(.A(new_n287), .B(new_n717), .C1(new_n707), .C2(new_n708), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n555), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n226), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n715), .A2(new_n722), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n719), .A2(new_n224), .A3(new_n514), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT100), .A2(KEYINPUT46), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT100), .A2(KEYINPUT46), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT101), .B1(new_n714), .B2(new_n552), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G36gat), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n714), .A2(KEYINPUT101), .A3(new_n552), .ZN(new_n730));
  OAI221_X1 g529(.A(new_n727), .B1(new_n725), .B2(new_n724), .C1(new_n729), .C2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n686), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n706), .A2(new_n732), .A3(new_n709), .A4(new_n713), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n688), .A2(new_n232), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n718), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n736), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n592), .A2(KEYINPUT103), .A3(new_n717), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT102), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT47), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n734), .A2(new_n740), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n742), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n744), .B2(new_n747), .ZN(G1330gat));
  OAI21_X1  g547(.A(new_n230), .B1(new_n718), .B2(new_n361), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n362), .A2(G50gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n714), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g551(.A1(new_n288), .A2(new_n648), .A3(new_n670), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n705), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n555), .B(KEYINPUT105), .Z(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n514), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT49), .B(G64gat), .Z(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(G1333gat));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n688), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n630), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n754), .A2(G71gat), .A3(new_n732), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n362), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n287), .A2(new_n711), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n670), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT107), .Z(new_n774));
  NAND2_X1  g573(.A1(new_n710), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n555), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n586), .A2(new_n686), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n558), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n625), .A3(new_n772), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n778), .A2(KEYINPUT51), .A3(new_n625), .A4(new_n772), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n603), .A3(new_n720), .A4(new_n670), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n784), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n775), .B2(new_n552), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n783), .A2(new_n604), .A3(new_n514), .A4(new_n670), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1337gat));
  XNOR2_X1  g591(.A(KEYINPUT108), .B(G99gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n783), .A2(new_n688), .A3(new_n670), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n775), .A2(new_n686), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n361), .A2(G106gat), .A3(new_n671), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT112), .B1(new_n783), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n706), .A2(new_n362), .A3(new_n709), .A4(new_n774), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT109), .B(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n783), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n799), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n797), .B(KEYINPUT110), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n781), .B2(new_n782), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n800), .A2(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n809), .B2(new_n810), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n814), .ZN(G1339gat));
  NOR4_X1   g614(.A1(new_n287), .A2(new_n625), .A3(new_n647), .A4(new_n670), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n251), .B1(new_n278), .B2(new_n250), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n269), .A2(new_n250), .A3(new_n267), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n205), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n286), .A2(new_n670), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n658), .A2(new_n654), .A3(new_n659), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n666), .B1(new_n660), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n825), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n669), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n280), .B2(new_n286), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n817), .B1(new_n821), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n830), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n272), .A2(new_n206), .A3(new_n279), .ZN(new_n834));
  INV_X1    g633(.A(new_n207), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n282), .B2(new_n285), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n286), .A2(new_n670), .A3(new_n820), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n832), .A2(new_n624), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n624), .A2(new_n830), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n286), .A3(new_n820), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n816), .B1(new_n843), .B2(new_n647), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n755), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n550), .A2(new_n551), .A3(new_n514), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n288), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n844), .A2(new_n362), .A3(new_n689), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n555), .A2(new_n514), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n287), .A2(G113gat), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n849), .A2(G113gat), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n852), .B2(new_n671), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n671), .A2(G120gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT116), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n848), .B2(new_n859), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n852), .B2(new_n647), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n647), .A2(G127gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n848), .B2(new_n862), .ZN(G1342gat));
  OR3_X1    g662(.A1(new_n848), .A2(G134gat), .A3(new_n624), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n852), .B2(new_n624), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n732), .A2(new_n514), .A3(new_n361), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n846), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n288), .A2(G141gat), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT58), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n829), .A2(new_n669), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT55), .B1(new_n826), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n825), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n287), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n624), .B1(new_n879), .B2(new_n821), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n842), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n816), .B1(new_n881), .B2(new_n647), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n361), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n711), .B1(new_n840), .B2(new_n842), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n362), .B1(new_n887), .B2(new_n816), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n686), .A2(new_n851), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n889), .A2(new_n288), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n872), .B1(new_n873), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT118), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n888), .A2(new_n883), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n886), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n287), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n898), .A2(G141gat), .B1(new_n870), .B2(new_n871), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n893), .A2(new_n897), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n902), .B(G148gat), .C1(new_n903), .C2(new_n671), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n884), .B1(new_n887), .B2(new_n816), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT119), .B(new_n884), .C1(new_n887), .C2(new_n816), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n286), .A2(new_n820), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n841), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n910), .B2(new_n841), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n711), .B1(new_n880), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n362), .B1(new_n913), .B2(new_n816), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n883), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n670), .A3(new_n895), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G148gat), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT121), .B1(new_n918), .B2(KEYINPUT59), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n920), .B(new_n902), .C1(new_n917), .C2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n904), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G148gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n870), .A2(new_n923), .A3(new_n670), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1345gat));
  OAI21_X1  g724(.A(G155gat), .B1(new_n903), .B2(new_n647), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n870), .A2(new_n292), .A3(new_n711), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1346gat));
  NAND3_X1  g727(.A1(new_n870), .A2(new_n293), .A3(new_n625), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT122), .ZN(new_n930));
  OAI21_X1  g729(.A(G162gat), .B1(new_n903), .B2(new_n624), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n844), .A2(new_n720), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT123), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n936), .A2(new_n383), .A3(new_n385), .A4(new_n287), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n755), .A2(new_n552), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n850), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n288), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(new_n940), .ZN(G1348gat));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n384), .A3(new_n670), .ZN(new_n942));
  OAI21_X1  g741(.A(G176gat), .B1(new_n939), .B2(new_n671), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  AND4_X1   g743(.A1(new_n395), .A2(new_n933), .A3(new_n711), .A4(new_n934), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n939), .A2(new_n647), .B1(new_n445), .B2(new_n444), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n396), .A3(new_n625), .ZN(new_n954));
  OAI21_X1  g753(.A(G190gat), .B1(new_n939), .B2(new_n624), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  AND4_X1   g758(.A1(new_n514), .A2(new_n933), .A3(new_n362), .A4(new_n686), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n287), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n686), .A2(new_n938), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n905), .A2(new_n906), .B1(new_n914), .B2(new_n883), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n908), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n287), .A2(G197gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n960), .A2(new_n967), .A3(new_n670), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  AOI211_X1 g768(.A(new_n671), .B(new_n962), .C1(new_n963), .C2(new_n908), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n967), .B2(new_n970), .ZN(G1353gat));
  INV_X1    g770(.A(G211gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n960), .A2(new_n972), .A3(new_n711), .ZN(new_n973));
  OAI21_X1  g772(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n964), .B2(new_n711), .ZN(new_n975));
  NAND2_X1  g774(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g776(.A(new_n647), .B(new_n962), .C1(new_n963), .C2(new_n908), .ZN(new_n978));
  INV_X1    g777(.A(new_n976), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(new_n974), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT126), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n976), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n978), .B2(new_n974), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n973), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n985), .ZN(G1354gat));
  NAND2_X1  g785(.A1(new_n964), .A2(new_n625), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n624), .A2(G218gat), .ZN(new_n988));
  AOI22_X1  g787(.A1(new_n987), .A2(G218gat), .B1(new_n960), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


