

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n725), .ZN(n690) );
  NAND2_X1 U550 ( .A1(G8), .A2(n725), .ZN(n723) );
  AND2_X2 U551 ( .A1(n687), .A2(n686), .ZN(n689) );
  NOR2_X1 U552 ( .A1(n689), .A2(n979), .ZN(n688) );
  OR2_X4 U553 ( .A1(G164), .A2(n683), .ZN(n725) );
  XOR2_X2 U554 ( .A(KEYINPUT89), .B(n526), .Z(G164) );
  XNOR2_X2 U555 ( .A(n517), .B(KEYINPUT65), .ZN(n675) );
  INV_X1 U556 ( .A(KEYINPUT103), .ZN(n731) );
  XNOR2_X1 U557 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U558 ( .A1(n863), .A2(G138), .ZN(n516) );
  INV_X1 U559 ( .A(KEYINPUT17), .ZN(n514) );
  NOR2_X1 U560 ( .A1(G651), .A2(n607), .ZN(n636) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XNOR2_X2 U562 ( .A(n515), .B(n514), .ZN(n863) );
  XOR2_X1 U563 ( .A(n516), .B(KEYINPUT87), .Z(n519) );
  INV_X1 U564 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n521), .A2(G2104), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n675), .A2(G102), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U568 ( .A(n520), .B(KEYINPUT88), .ZN(n525) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n866) );
  NAND2_X1 U570 ( .A1(G114), .A2(n866), .ZN(n523) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n521), .ZN(n867) );
  NAND2_X1 U572 ( .A1(G126), .A2(n867), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n527) );
  XNOR2_X1 U576 ( .A(n527), .B(KEYINPUT64), .ZN(n639) );
  NAND2_X1 U577 ( .A1(G89), .A2(n639), .ZN(n528) );
  XNOR2_X1 U578 ( .A(n528), .B(KEYINPUT4), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n607) );
  INV_X1 U580 ( .A(G651), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n607), .A2(n532), .ZN(n642) );
  NAND2_X1 U582 ( .A1(G76), .A2(n642), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U584 ( .A(KEYINPUT5), .B(n531), .ZN(n539) );
  NOR2_X1 U585 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n533), .Z(n638) );
  NAND2_X1 U587 ( .A1(G63), .A2(n638), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G51), .A2(n636), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT74), .B(KEYINPUT6), .Z(n536) );
  XNOR2_X1 U591 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U593 ( .A(KEYINPUT7), .B(n540), .ZN(G168) );
  XOR2_X1 U594 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U595 ( .A1(n642), .A2(G78), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G91), .A2(n639), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U598 ( .A(KEYINPUT67), .B(n543), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G65), .A2(n638), .ZN(n544) );
  XOR2_X1 U600 ( .A(KEYINPUT68), .B(n544), .Z(n547) );
  NAND2_X1 U601 ( .A1(G53), .A2(n636), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT69), .B(n545), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(G299) );
  XOR2_X1 U605 ( .A(G2438), .B(G2454), .Z(n551) );
  XNOR2_X1 U606 ( .A(G2435), .B(G2430), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U608 ( .A(n552), .B(G2427), .Z(n554) );
  XNOR2_X1 U609 ( .A(G1348), .B(G1341), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U611 ( .A(G2443), .B(G2446), .Z(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT106), .B(G2451), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U614 ( .A(n558), .B(n557), .Z(n559) );
  AND2_X1 U615 ( .A1(G14), .A2(n559), .ZN(G401) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U617 ( .A1(G135), .A2(n863), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G111), .A2(n866), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n867), .A2(G123), .ZN(n562) );
  XOR2_X1 U621 ( .A(KEYINPUT18), .B(n562), .Z(n563) );
  NOR2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n675), .A2(G99), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n921) );
  XNOR2_X1 U625 ( .A(G2096), .B(n921), .ZN(n567) );
  OR2_X1 U626 ( .A1(G2100), .A2(n567), .ZN(G156) );
  NAND2_X1 U627 ( .A1(n642), .A2(G77), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G90), .A2(n639), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n570), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G64), .A2(n638), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G52), .A2(n636), .ZN(n571) );
  AND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G301) );
  INV_X1 U635 ( .A(G301), .ZN(G171) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n830) );
  NAND2_X1 U639 ( .A1(n830), .A2(G567), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n638), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U643 ( .A1(G81), .A2(n639), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G68), .A2(n642), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n636), .A2(G43), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n976) );
  INV_X1 U651 ( .A(G860), .ZN(n598) );
  OR2_X1 U652 ( .A1(n976), .A2(n598), .ZN(G153) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U654 ( .A1(G79), .A2(n642), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G54), .A2(n636), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G92), .A2(n639), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G66), .A2(n638), .ZN(n588) );
  XNOR2_X1 U659 ( .A(KEYINPUT73), .B(n588), .ZN(n589) );
  NOR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT15), .ZN(n979) );
  OR2_X1 U663 ( .A1(n979), .A2(G868), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G284) );
  INV_X1 U665 ( .A(G868), .ZN(n657) );
  NOR2_X1 U666 ( .A1(G286), .A2(n657), .ZN(n597) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n979), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT75), .B(n601), .Z(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n976), .ZN(n602) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n602), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G868), .A2(n979), .ZN(n603) );
  NOR2_X1 U676 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G74), .A2(G651), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT82), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G49), .A2(n636), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G87), .A2(n607), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n638), .A2(n610), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT83), .B(n613), .Z(G288) );
  NAND2_X1 U686 ( .A1(G62), .A2(n638), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G88), .A2(n639), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G75), .A2(n642), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT85), .B(n616), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n636), .A2(G50), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G303) );
  INV_X1 U694 ( .A(G303), .ZN(G166) );
  NAND2_X1 U695 ( .A1(G60), .A2(n638), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G47), .A2(n636), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U698 ( .A(KEYINPUT66), .B(n623), .Z(n627) );
  NAND2_X1 U699 ( .A1(n639), .A2(G85), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n642), .A2(G72), .ZN(n624) );
  AND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(G290) );
  XOR2_X1 U703 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n629) );
  NAND2_X1 U704 ( .A1(G73), .A2(n642), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n629), .B(n628), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G61), .A2(n638), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G86), .A2(n639), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(G48), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U712 ( .A1(G55), .A2(n636), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT80), .ZN(n647) );
  NAND2_X1 U714 ( .A1(G67), .A2(n638), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G93), .A2(n639), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U717 ( .A1(G80), .A2(n642), .ZN(n643) );
  XNOR2_X1 U718 ( .A(KEYINPUT79), .B(n643), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT81), .B(n648), .Z(n841) );
  XNOR2_X1 U722 ( .A(G166), .B(KEYINPUT19), .ZN(n650) );
  INV_X1 U723 ( .A(G299), .ZN(n969) );
  XNOR2_X1 U724 ( .A(G290), .B(n969), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U726 ( .A(n651), .B(G305), .Z(n652) );
  XNOR2_X1 U727 ( .A(G288), .B(n652), .ZN(n653) );
  XOR2_X1 U728 ( .A(n841), .B(n653), .Z(n885) );
  XNOR2_X1 U729 ( .A(n976), .B(KEYINPUT77), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n979), .A2(G559), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n838) );
  XNOR2_X1 U732 ( .A(n885), .B(n838), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n656), .A2(G868), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n657), .A2(n841), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XOR2_X1 U741 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U743 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U744 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NAND2_X1 U745 ( .A1(G120), .A2(G69), .ZN(n664) );
  NOR2_X1 U746 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U747 ( .A1(G108), .A2(n665), .ZN(n836) );
  NAND2_X1 U748 ( .A1(n836), .A2(G567), .ZN(n670) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U751 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G96), .A2(n668), .ZN(n835) );
  NAND2_X1 U753 ( .A1(n835), .A2(G2106), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n842) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n671) );
  XNOR2_X1 U756 ( .A(KEYINPUT86), .B(n671), .ZN(n672) );
  NOR2_X1 U757 ( .A1(n842), .A2(n672), .ZN(n834) );
  NAND2_X1 U758 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(G113), .A2(n866), .ZN(n674) );
  NAND2_X1 U760 ( .A1(G125), .A2(n867), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G101), .A2(n675), .ZN(n676) );
  XOR2_X1 U763 ( .A(KEYINPUT23), .B(n676), .Z(n678) );
  NAND2_X1 U764 ( .A1(n863), .A2(G137), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U766 ( .A1(n680), .A2(n679), .ZN(G160) );
  INV_X1 U767 ( .A(G1384), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n762) );
  INV_X1 U769 ( .A(n762), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n690), .A2(G1996), .ZN(n684) );
  XNOR2_X1 U772 ( .A(n684), .B(KEYINPUT26), .ZN(n687) );
  AND2_X1 U773 ( .A1(n725), .A2(G1341), .ZN(n685) );
  NOR2_X1 U774 ( .A1(n685), .A2(n976), .ZN(n686) );
  XOR2_X1 U775 ( .A(n688), .B(KEYINPUT98), .Z(n696) );
  NAND2_X1 U776 ( .A1(n689), .A2(n979), .ZN(n694) );
  NOR2_X1 U777 ( .A1(G2067), .A2(n725), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n690), .A2(G1348), .ZN(n691) );
  NOR2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n696), .A2(n695), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n690), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U783 ( .A(n697), .B(KEYINPUT27), .ZN(n699) );
  INV_X1 U784 ( .A(G1956), .ZN(n994) );
  NOR2_X1 U785 ( .A1(n994), .A2(n690), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U787 ( .A1(n969), .A2(n702), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U789 ( .A1(n969), .A2(n702), .ZN(n704) );
  XNOR2_X1 U790 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n703) );
  XNOR2_X1 U791 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U793 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n707) );
  XNOR2_X1 U794 ( .A(n708), .B(n707), .ZN(n712) );
  XOR2_X1 U795 ( .A(G1961), .B(KEYINPUT96), .Z(n993) );
  NAND2_X1 U796 ( .A1(n993), .A2(n725), .ZN(n710) );
  XNOR2_X1 U797 ( .A(KEYINPUT25), .B(G2078), .ZN(n945) );
  NAND2_X1 U798 ( .A1(n690), .A2(n945), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U800 ( .A1(n716), .A2(G171), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n722) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n725), .ZN(n735) );
  NOR2_X1 U803 ( .A1(n723), .A2(G1966), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n735), .A2(n739), .ZN(n713) );
  NAND2_X1 U805 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n714), .B(KEYINPUT30), .ZN(n715) );
  NOR2_X1 U807 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U808 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U810 ( .A(KEYINPUT100), .B(n719), .Z(n720) );
  XNOR2_X1 U811 ( .A(KEYINPUT31), .B(n720), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n737), .A2(G286), .ZN(n730) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n723), .ZN(n724) );
  XNOR2_X1 U815 ( .A(n724), .B(KEYINPUT102), .ZN(n727) );
  NOR2_X1 U816 ( .A1(n725), .A2(G2090), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U818 ( .A1(n728), .A2(G303), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT32), .ZN(n796) );
  NAND2_X1 U822 ( .A1(G8), .A2(n735), .ZN(n736) );
  XOR2_X1 U823 ( .A(KEYINPUT95), .B(n736), .Z(n743) );
  INV_X1 U824 ( .A(KEYINPUT101), .ZN(n741) );
  INV_X1 U825 ( .A(n737), .ZN(n738) );
  NOR2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n789) );
  NOR2_X1 U829 ( .A1(G1981), .A2(G305), .ZN(n744) );
  XOR2_X1 U830 ( .A(n744), .B(KEYINPUT24), .Z(n745) );
  NOR2_X1 U831 ( .A1(n723), .A2(n745), .ZN(n782) );
  OR2_X1 U832 ( .A1(n782), .A2(n723), .ZN(n778) );
  NAND2_X1 U833 ( .A1(G107), .A2(n866), .ZN(n747) );
  NAND2_X1 U834 ( .A1(G119), .A2(n867), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G95), .A2(n675), .ZN(n748) );
  XNOR2_X1 U837 ( .A(KEYINPUT93), .B(n748), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n863), .A2(G131), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n876) );
  AND2_X1 U841 ( .A1(n876), .A2(G1991), .ZN(n761) );
  NAND2_X1 U842 ( .A1(G117), .A2(n866), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G129), .A2(n867), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n675), .A2(G105), .ZN(n755) );
  XOR2_X1 U846 ( .A(KEYINPUT38), .B(n755), .Z(n756) );
  NOR2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n863), .A2(G141), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n878) );
  AND2_X1 U850 ( .A1(n878), .A2(G1996), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n926) );
  NOR2_X1 U852 ( .A1(G164), .A2(G1384), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n825) );
  INV_X1 U854 ( .A(n825), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n926), .A2(n764), .ZN(n817) );
  INV_X1 U856 ( .A(n817), .ZN(n776) );
  NAND2_X1 U857 ( .A1(G140), .A2(n863), .ZN(n766) );
  NAND2_X1 U858 ( .A1(G104), .A2(n675), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n767), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G116), .A2(n866), .ZN(n769) );
  NAND2_X1 U862 ( .A1(G128), .A2(n867), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U864 ( .A(n770), .B(KEYINPUT35), .Z(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n773), .Z(n774) );
  XOR2_X1 U867 ( .A(KEYINPUT91), .B(n774), .Z(n860) );
  XOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .Z(n822) );
  AND2_X1 U869 ( .A1(n860), .A2(n822), .ZN(n775) );
  XNOR2_X1 U870 ( .A(n775), .B(KEYINPUT92), .ZN(n935) );
  NAND2_X1 U871 ( .A1(n825), .A2(n935), .ZN(n820) );
  NAND2_X1 U872 ( .A1(n776), .A2(n820), .ZN(n777) );
  XOR2_X1 U873 ( .A(n777), .B(KEYINPUT94), .Z(n790) );
  NAND2_X1 U874 ( .A1(n778), .A2(n790), .ZN(n786) );
  INV_X1 U875 ( .A(n786), .ZN(n779) );
  AND2_X1 U876 ( .A1(n789), .A2(n779), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n796), .A2(n780), .ZN(n788) );
  NOR2_X1 U878 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U879 ( .A1(G8), .A2(n781), .ZN(n784) );
  INV_X1 U880 ( .A(n782), .ZN(n783) );
  AND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n810) );
  NAND2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U885 ( .A1(n789), .A2(n974), .ZN(n794) );
  XOR2_X1 U886 ( .A(G1981), .B(G305), .Z(n984) );
  AND2_X1 U887 ( .A1(n984), .A2(n790), .ZN(n797) );
  NOR2_X1 U888 ( .A1(G1976), .A2(G288), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n799), .A2(KEYINPUT33), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n791), .A2(n723), .ZN(n804) );
  INV_X1 U891 ( .A(n804), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n797), .A2(n792), .ZN(n793) );
  NOR2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n808) );
  INV_X1 U895 ( .A(n797), .ZN(n806) );
  INV_X1 U896 ( .A(n974), .ZN(n800) );
  NOR2_X1 U897 ( .A1(G1971), .A2(G303), .ZN(n798) );
  NOR2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n983) );
  OR2_X1 U899 ( .A1(n800), .A2(n983), .ZN(n801) );
  NOR2_X1 U900 ( .A1(n723), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n802), .A2(KEYINPUT33), .ZN(n803) );
  OR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X2 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U906 ( .A(n811), .B(KEYINPUT104), .ZN(n814) );
  XNOR2_X1 U907 ( .A(KEYINPUT90), .B(G1986), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(G290), .ZN(n973) );
  NAND2_X1 U909 ( .A1(n973), .A2(n825), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n828) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n878), .ZN(n928) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n876), .ZN(n924) );
  NOR2_X1 U914 ( .A1(n815), .A2(n924), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n928), .A2(n818), .ZN(n819) );
  XNOR2_X1 U917 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n860), .A2(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT105), .ZN(n932) );
  NAND2_X1 U921 ( .A1(n824), .A2(n932), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(n830), .A2(G2106), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT107), .B(n831), .Z(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U928 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U931 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NOR2_X1 U936 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n837), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U938 ( .A(G261), .ZN(G325) );
  XOR2_X1 U939 ( .A(KEYINPUT78), .B(n838), .Z(n839) );
  NOR2_X1 U940 ( .A1(G860), .A2(n839), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(G145) );
  INV_X1 U942 ( .A(n842), .ZN(G319) );
  NAND2_X1 U943 ( .A1(G124), .A2(n867), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n843), .B(KEYINPUT112), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G112), .A2(n866), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U948 ( .A1(G136), .A2(n863), .ZN(n848) );
  NAND2_X1 U949 ( .A1(G100), .A2(n675), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U951 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G142), .A2(n863), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G106), .A2(n675), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT45), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G130), .A2(n867), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G118), .A2(n866), .ZN(n856) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(n856), .ZN(n857) );
  NOR2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n921), .B(n859), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n860), .B(G162), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n883) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n875) );
  NAND2_X1 U965 ( .A1(G139), .A2(n863), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G103), .A2(n675), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G115), .A2(n866), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G127), .A2(n867), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(n871), .ZN(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n915) );
  XNOR2_X1 U974 ( .A(n915), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n880) );
  XOR2_X1 U977 ( .A(G160), .B(n878), .Z(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U981 ( .A1(G37), .A2(n884), .ZN(G395) );
  XOR2_X1 U982 ( .A(n885), .B(G286), .Z(n887) );
  XNOR2_X1 U983 ( .A(G171), .B(n979), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(n888), .B(n976), .Z(n889) );
  NOR2_X1 U986 ( .A1(G37), .A2(n889), .ZN(G397) );
  XOR2_X1 U987 ( .A(KEYINPUT110), .B(G1981), .Z(n891) );
  XNOR2_X1 U988 ( .A(G1966), .B(G1956), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n892), .B(G2474), .Z(n894) );
  XNOR2_X1 U991 ( .A(G1996), .B(G1991), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U993 ( .A(G1976), .B(G1971), .Z(n896) );
  XNOR2_X1 U994 ( .A(G1986), .B(G1961), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n900) );
  XNOR2_X1 U997 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(G229) );
  XOR2_X1 U999 ( .A(G2100), .B(G2096), .Z(n902) );
  XNOR2_X1 U1000 ( .A(KEYINPUT42), .B(G2678), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1002 ( .A(KEYINPUT43), .B(G2090), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G2072), .B(G2067), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1006 ( .A(G2084), .B(G2078), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(G227) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT116), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n912) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1016 ( .A(G2072), .B(n915), .Z(n917) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(n918), .B(KEYINPUT50), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n920), .B(n919), .ZN(n938) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n931) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n929), .B(KEYINPUT51), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n965) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n965), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n941), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1038 ( .A(G2072), .B(G33), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G26), .B(G2067), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1041 ( .A(KEYINPUT122), .B(n944), .Z(n950) );
  XOR2_X1 U1042 ( .A(n945), .B(G27), .Z(n947) );
  XNOR2_X1 U1043 ( .A(G32), .B(G1996), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT123), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1047 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1048 ( .A1(n951), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(KEYINPUT121), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(KEYINPUT53), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT124), .B(n956), .ZN(n963) );
  XOR2_X1 U1053 ( .A(KEYINPUT125), .B(G34), .Z(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(KEYINPUT126), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n958), .B(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G2090), .B(G35), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1061 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n968), .ZN(n1021) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1065 ( .A(n969), .B(G1956), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n976), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n990) );
  XOR2_X1 U1072 ( .A(G1348), .B(n979), .Z(n981) );
  XOR2_X1 U1073 ( .A(G171), .B(G1961), .Z(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n1019) );
  INV_X1 U1082 ( .A(G16), .ZN(n1017) );
  XNOR2_X1 U1083 ( .A(n993), .B(G5), .ZN(n1007) );
  XNOR2_X1 U1084 ( .A(G20), .B(n994), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1090 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n1002) );
  XOR2_X1 U1093 ( .A(n1003), .B(n1002), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G21), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(G1986), .B(G24), .Z(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

