//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G113gat), .B2(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G113gat), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n205), .A3(new_n207), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(new_n210), .A3(new_n204), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT68), .B1(new_n212), .B2(new_n217), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G183gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n222), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G183gat), .B(G190gat), .ZN(new_n232));
  OAI211_X1 g031(.A(KEYINPUT64), .B(new_n229), .C1(new_n232), .C2(new_n223), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT23), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n229), .B1(new_n232), .B2(new_n223), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n246), .A2(new_n239), .A3(new_n243), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n226), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n250), .A2(KEYINPUT66), .A3(KEYINPUT28), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n252));
  AND2_X1   g051(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n253));
  AOI211_X1 g052(.A(new_n252), .B(new_n253), .C1(new_n249), .C2(new_n226), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n234), .A2(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n236), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n234), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n251), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n221), .B1(new_n248), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n243), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n265));
  INV_X1    g064(.A(new_n247), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n220), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n218), .ZN(new_n269));
  INV_X1    g068(.A(new_n259), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n260), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT33), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n283), .B2(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT34), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n262), .B1(new_n260), .B2(new_n271), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT72), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n247), .B1(new_n263), .B2(KEYINPUT65), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n259), .B(new_n221), .C1(new_n294), .C2(new_n265), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n269), .B1(new_n267), .B2(new_n270), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n261), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n297), .B2(KEYINPUT71), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT34), .B1(new_n297), .B2(new_n293), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n288), .B(new_n292), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n290), .B2(new_n291), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n289), .B1(new_n290), .B2(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n288), .B1(new_n304), .B2(new_n292), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n287), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(new_n286), .A3(new_n282), .A4(new_n300), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n309), .A3(KEYINPUT74), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT36), .ZN(new_n311));
  INV_X1    g110(.A(new_n287), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n312), .A2(new_n313), .A3(new_n308), .A4(new_n300), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n306), .A2(new_n309), .A3(KEYINPUT36), .ZN(new_n316));
  XNOR2_X1  g115(.A(G1gat), .B(G29gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT0), .ZN(new_n318));
  XNOR2_X1  g117(.A(G57gat), .B(G85gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(G141gat), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n325), .A2(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT81), .B(G155gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n333), .B2(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G148gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G141gat), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n327), .A2(new_n341), .B1(KEYINPUT2), .B2(new_n331), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT78), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT78), .B1(new_n328), .B2(new_n329), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n331), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT79), .B(new_n331), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n212), .A2(new_n217), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n339), .B2(new_n349), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n322), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n332), .A2(new_n337), .A3(new_n334), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n337), .B1(new_n332), .B2(new_n334), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g157(.A(new_n350), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n349), .B(new_n360), .C1(new_n355), .C2(new_n356), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n321), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n221), .A2(new_n339), .A3(KEYINPUT4), .A4(new_n349), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n352), .B2(KEYINPUT4), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT5), .B(new_n354), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n357), .B2(new_n269), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n349), .A4(new_n350), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n321), .A4(new_n362), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n320), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT6), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n372), .A3(new_n320), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT83), .ZN(new_n378));
  INV_X1    g177(.A(new_n373), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n377), .A2(KEYINPUT83), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386));
  AND2_X1   g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n385), .A2(KEYINPUT22), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G211gat), .B(G218gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n267), .A2(new_n270), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(KEYINPUT75), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT76), .B1(new_n248), .B2(new_n259), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n267), .A2(new_n397), .A3(new_n270), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n391), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n394), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n390), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(KEYINPUT77), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n398), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n397), .B1(new_n267), .B2(new_n270), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n393), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n391), .A4(new_n395), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT30), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n410), .B1(new_n406), .B2(new_n416), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT30), .B(new_n410), .C1(new_n406), .C2(new_n416), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n382), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n391), .B1(new_n361), .B2(new_n403), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n360), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n357), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n424), .A2(new_n426), .A3(new_n423), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n428), .A2(G22gat), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(G22gat), .B1(new_n428), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n428), .A2(new_n429), .A3(G22gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(KEYINPUT84), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n315), .A2(new_n316), .B1(new_n422), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT39), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n361), .A2(new_n359), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n360), .B1(new_n339), .B2(new_n349), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n368), .B(new_n369), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n446), .A2(new_n447), .A3(new_n322), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n446), .B2(new_n322), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n322), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n446), .A2(new_n447), .A3(new_n322), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n352), .A2(new_n353), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n454), .B2(new_n321), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n456), .A3(new_n320), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n379), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(KEYINPUT86), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n450), .A2(new_n456), .A3(new_n461), .A4(new_n320), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n421), .ZN(new_n466));
  INV_X1    g265(.A(new_n419), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n417), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n460), .A2(KEYINPUT87), .A3(new_n458), .A4(new_n462), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT37), .B1(new_n406), .B2(new_n416), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n402), .A2(new_n404), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n391), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n414), .A2(new_n390), .A3(new_n395), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT38), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n410), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n374), .B1(new_n377), .B2(new_n373), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n419), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n406), .A2(KEYINPUT37), .A3(new_n416), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n481), .A2(new_n471), .A3(new_n409), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT38), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n478), .B(new_n480), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n470), .A2(new_n440), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n442), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n306), .A2(new_n309), .A3(new_n440), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n422), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n310), .A2(new_n314), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n466), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n440), .A2(new_n491), .A3(new_n479), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G57gat), .B(G64gat), .Z(new_n496));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497));
  INV_X1    g296(.A(G71gat), .ZN(new_n498));
  INV_X1    g297(.A(G78gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(new_n203), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(G1gat), .B2(new_n509), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G8gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n501), .B(new_n502), .Z(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(KEYINPUT21), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n508), .B(new_n515), .Z(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n328), .ZN(new_n518));
  XNOR2_X1  g317(.A(G183gat), .B(G211gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n518), .B(new_n519), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n508), .B(new_n515), .ZN(new_n522));
  INV_X1    g321(.A(new_n520), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G230gat), .ZN(new_n526));
  INV_X1    g325(.A(G233gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g328(.A(G85gat), .ZN(new_n530));
  INV_X1    g329(.A(G92gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  AOI22_X1  g334(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n530), .B2(new_n531), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G99gat), .B(G106gat), .Z(new_n538));
  OR2_X1    g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT98), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n543), .A3(new_n503), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n514), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT100), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT10), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT100), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n539), .A2(new_n514), .A3(new_n548), .A4(new_n540), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT10), .A3(new_n514), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n528), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n528), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(G176gat), .B(G204gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT96), .ZN(new_n569));
  XOR2_X1   g368(.A(G134gat), .B(G162gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G43gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G50gat), .ZN(new_n573));
  INV_X1    g372(.A(G50gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(G43gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n576));
  OR3_X1    g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n573), .B2(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT15), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(new_n573), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n572), .A3(G50gat), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT15), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OR3_X1    g383(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT14), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(KEYINPUT14), .ZN(new_n588));
  INV_X1    g387(.A(G29gat), .ZN(new_n589));
  INV_X1    g388(.A(G36gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT90), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT90), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n587), .A2(new_n588), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n579), .B1(new_n584), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n579), .B2(new_n593), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT92), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n551), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(KEYINPUT17), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT93), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n596), .A2(new_n551), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n571), .B1(new_n605), .B2(KEYINPUT99), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(new_n604), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n601), .B2(new_n602), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR4_X1   g410(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT99), .A4(new_n571), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n525), .B(new_n566), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT94), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n596), .A2(new_n513), .ZN(new_n616));
  INV_X1    g415(.A(new_n513), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n595), .B(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n619), .B2(KEYINPUT17), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n599), .B(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n615), .B(new_n616), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n600), .B(new_n617), .C1(KEYINPUT17), .C2(new_n619), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n626), .A2(KEYINPUT18), .A3(new_n615), .A4(new_n616), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n596), .B2(new_n513), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(KEYINPUT95), .A3(new_n617), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n616), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n615), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G197gat), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT11), .B(G169gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n627), .A3(new_n641), .A4(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n613), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n495), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n382), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  INV_X1    g450(.A(new_n490), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT16), .B(G8gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(G8gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(KEYINPUT42), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(G1325gat));
  NAND2_X1  g458(.A1(new_n315), .A2(new_n316), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n489), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n646), .B2(new_n663), .ZN(G1326gat));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n440), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n611), .A2(new_n612), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n495), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n644), .A2(new_n525), .A3(new_n565), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n589), .A3(new_n648), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n495), .A2(KEYINPUT44), .A3(new_n668), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n442), .A2(new_n485), .B1(new_n488), .B2(new_n493), .ZN(new_n677));
  INV_X1    g476(.A(new_n668), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n382), .A3(new_n671), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n674), .B1(new_n589), .B2(new_n681), .ZN(G1328gat));
  NAND3_X1  g481(.A1(new_n672), .A2(new_n590), .A3(new_n652), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT46), .Z(new_n684));
  NOR2_X1   g483(.A1(new_n680), .A2(new_n671), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n652), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G36gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(new_n660), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n685), .A2(G43gat), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n672), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n572), .B1(new_n693), .B2(new_n662), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g495(.A1(new_n672), .A2(new_n574), .A3(new_n441), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n440), .A3(new_n671), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(new_n574), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT48), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n699), .B(new_n701), .ZN(G1331gat));
  AND2_X1   g501(.A1(new_n521), .A2(new_n524), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n704), .A2(new_n571), .B1(new_n607), .B2(new_n609), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n606), .A2(new_n610), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n495), .A2(new_n644), .A3(new_n707), .A4(new_n565), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n648), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT104), .B(G57gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n652), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT49), .B(G64gat), .Z(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(G1333gat));
  AOI21_X1  g514(.A(new_n498), .B1(new_n708), .B2(new_n691), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n662), .A2(G71gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n708), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n708), .A2(new_n441), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g520(.A(new_n678), .B1(new_n486), .B2(new_n494), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n643), .A2(new_n525), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT51), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  INV_X1    g524(.A(new_n723), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n677), .A2(new_n725), .A3(new_n678), .A4(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n566), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n530), .A3(new_n648), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n726), .A2(new_n566), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n675), .A2(new_n679), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n675), .A2(new_n679), .A3(KEYINPUT105), .A4(new_n731), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(new_n648), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n736), .B2(new_n530), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT106), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n652), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G92gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n677), .A2(new_n678), .A3(new_n726), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n725), .B1(new_n741), .B2(KEYINPUT107), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(KEYINPUT51), .C1(new_n669), .C2(new_n726), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n490), .A2(G92gat), .A3(new_n566), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(KEYINPUT108), .A3(KEYINPUT52), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n739), .A2(G92gat), .B1(new_n745), .B2(new_n746), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n746), .B1(new_n724), .B2(new_n727), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT109), .B(new_n746), .C1(new_n724), .C2(new_n727), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n675), .A2(new_n679), .A3(new_n652), .A4(new_n731), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n531), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n760), .B2(new_n759), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT111), .B1(new_n758), .B2(new_n762), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n749), .B(new_n753), .C1(new_n763), .C2(new_n764), .ZN(G1337gat));
  INV_X1    g564(.A(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n729), .A2(new_n766), .A3(new_n489), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n734), .A2(new_n691), .A3(new_n735), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n766), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1338gat));
  NOR3_X1   g570(.A1(new_n566), .A2(new_n440), .A3(G106gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n742), .A2(new_n744), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n734), .A2(new_n441), .A3(new_n735), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G106gat), .B1(new_n732), .B2(new_n440), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n772), .B1(new_n724), .B2(new_n727), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n652), .A2(new_n382), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n615), .B1(new_n626), .B2(new_n616), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n631), .A2(new_n632), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n638), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n642), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n565), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n550), .A2(new_n528), .A3(new_n552), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n553), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n560), .B1(new_n553), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT54), .B(new_n528), .C1(new_n550), .C2(new_n552), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(new_n560), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n795), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n791), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n799), .B1(new_n798), .B2(new_n560), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n794), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n562), .B1(new_n806), .B2(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n643), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n790), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n678), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n803), .A2(new_n807), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n813), .A2(new_n668), .A3(new_n789), .A4(new_n809), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n703), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n707), .A2(KEYINPUT114), .A3(new_n644), .A4(new_n566), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n613), .B2(new_n643), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n487), .B(new_n785), .C1(new_n816), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n643), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n441), .B1(new_n816), .B2(new_n821), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(new_n489), .A3(new_n784), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n644), .A2(new_n213), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(G120gat), .B1(new_n822), .B2(new_n565), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n566), .A2(new_n214), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1341gat));
  NAND3_X1  g629(.A1(new_n825), .A2(G127gat), .A3(new_n525), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n833));
  AOI21_X1  g632(.A(G127gat), .B1(new_n822), .B2(new_n525), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n822), .A2(new_n836), .A3(new_n668), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n825), .B2(new_n668), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(KEYINPUT56), .B2(new_n837), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n801), .A2(new_n802), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n643), .A2(new_n809), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n790), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n678), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n525), .B1(new_n845), .B2(new_n814), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n441), .B1(new_n846), .B2(new_n820), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n525), .B1(new_n812), .B2(new_n814), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n849), .B(new_n441), .C1(new_n850), .C2(new_n820), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n785), .A2(new_n691), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n848), .A2(new_n851), .A3(new_n643), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n326), .B1(new_n853), .B2(KEYINPUT120), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(KEYINPUT120), .B2(new_n853), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n816), .A2(new_n821), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n441), .A2(new_n857), .A3(new_n660), .A4(new_n784), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n326), .A3(new_n643), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(G141gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n853), .A2(new_n863), .A3(G141gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n864), .A3(new_n859), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT58), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n865), .B2(KEYINPUT58), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n323), .A2(new_n324), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n858), .A2(new_n871), .A3(new_n565), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n613), .A2(new_n643), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n849), .B(new_n441), .C1(new_n846), .C2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n440), .B1(new_n816), .B2(new_n821), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n849), .ZN(new_n878));
  OR4_X1    g677(.A1(new_n691), .A2(new_n878), .A3(new_n566), .A4(new_n785), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n871), .C1(new_n881), .C2(new_n565), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n880), .B2(new_n882), .ZN(G1345gat));
  NAND3_X1  g682(.A1(new_n858), .A2(new_n333), .A3(new_n525), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n881), .A2(new_n525), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n333), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n858), .B2(new_n668), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n678), .A2(new_n329), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n881), .B2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n490), .A2(new_n648), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n487), .B(new_n891), .C1(new_n816), .C2(new_n821), .ZN(new_n892));
  INV_X1    g691(.A(G169gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n643), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT122), .Z(new_n895));
  NOR2_X1   g694(.A1(new_n891), .A2(new_n662), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n824), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n644), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1348gat));
  NAND4_X1  g698(.A1(new_n824), .A2(G176gat), .A3(new_n565), .A4(new_n896), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  AOI21_X1  g702(.A(G176gat), .B1(new_n892), .B2(new_n565), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G1349gat));
  OAI21_X1  g704(.A(G183gat), .B1(new_n897), .B2(new_n703), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n892), .A2(new_n249), .A3(new_n525), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n226), .A3(new_n668), .ZN(new_n910));
  OAI21_X1  g709(.A(G190gat), .B1(new_n897), .B2(new_n678), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1351gat));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n878), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT124), .B(new_n876), .C1(new_n877), .C2(new_n849), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n691), .A2(new_n891), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G197gat), .B1(new_n919), .B2(new_n644), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n877), .A2(new_n918), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n921), .A2(G197gat), .A3(new_n644), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1352gat));
  OAI21_X1  g726(.A(G204gat), .B1(new_n919), .B2(new_n566), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n921), .A2(G204gat), .A3(new_n566), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  NAND4_X1  g730(.A1(new_n877), .A2(new_n383), .A3(new_n525), .A4(new_n918), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n691), .A2(new_n703), .A3(new_n891), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G211gat), .B1(new_n878), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(new_n384), .B1(new_n921), .B2(new_n678), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n668), .A2(G218gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n919), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


