//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT77), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n206), .A2(new_n209), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g021(.A(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n208), .A2(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n221), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n214), .B2(new_n220), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT78), .A3(new_n222), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT29), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT72), .B(G211gat), .ZN(new_n237));
  INV_X1    g036(.A(G218gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT73), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n240), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n203), .B1(new_n235), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n233), .B2(new_n222), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n219), .B1(new_n211), .B2(new_n213), .ZN(new_n252));
  NOR4_X1   g051(.A1(new_n252), .A2(new_n231), .A3(KEYINPUT3), .A4(new_n228), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT84), .A3(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n222), .B1(new_n247), .B2(KEYINPUT29), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n221), .A2(new_n229), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n256), .B(KEYINPUT82), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n232), .A2(new_n234), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n248), .B1(new_n262), .B2(new_n250), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT83), .B1(new_n239), .B2(new_n240), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n242), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n244), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n264), .B2(new_n242), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n233), .B1(new_n269), .B2(new_n222), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n261), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n202), .B1(new_n260), .B2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n260), .A2(new_n202), .A3(new_n271), .ZN(new_n274));
  XOR2_X1   g073(.A(G78gat), .B(G106gat), .Z(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT31), .B(G50gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n271), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G22gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n202), .A3(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT85), .B1(new_n284), .B2(new_n277), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT85), .B(new_n277), .C1(new_n274), .C2(new_n272), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n280), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n293));
  AND3_X1   g092(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT24), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n293), .B(KEYINPUT65), .C1(new_n294), .C2(new_n295), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(KEYINPUT25), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n298), .A2(new_n308), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n293), .B(new_n311), .C1(new_n294), .C2(new_n295), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n304), .A2(new_n306), .B1(new_n300), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n300), .A2(KEYINPUT27), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G183gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n299), .A2(new_n319), .A3(new_n321), .A4(new_n301), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n301), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT27), .B(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n323), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n303), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n294), .A2(new_n295), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n313), .A2(new_n318), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n349), .ZN(new_n351));
  XNOR2_X1  g150(.A(G113gat), .B(G120gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(KEYINPUT1), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n313), .A2(new_n318), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n338), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n357), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n290), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n360), .B(KEYINPUT32), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n360), .B2(KEYINPUT32), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n358), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n354), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n339), .A2(new_n355), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n289), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT33), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT68), .B1(new_n360), .B2(new_n361), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n366), .B(new_n367), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n371), .B2(KEYINPUT33), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n360), .A2(KEYINPUT68), .A3(new_n361), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n366), .B1(new_n379), .B2(new_n367), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n365), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n369), .A2(new_n289), .A3(new_n370), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT34), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n289), .B2(KEYINPUT70), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n384), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n379), .A2(new_n367), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT69), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n375), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n365), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n288), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n355), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n251), .B2(new_n253), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n221), .A2(new_n229), .A3(new_n355), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT4), .B1(new_n233), .B2(new_n355), .ZN(new_n412));
  NOR4_X1   g211(.A1(new_n252), .A2(new_n354), .A3(new_n408), .A4(new_n228), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT79), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n402), .B(new_n405), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n354), .B1(new_n252), .B2(new_n228), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n404), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n354), .B1(new_n233), .B2(new_n222), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n232), .B2(new_n234), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n409), .A2(new_n410), .A3(new_n403), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n415), .B2(new_n423), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n400), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n423), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n429), .A4(new_n428), .ZN(new_n436));
  INV_X1    g235(.A(new_n429), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n368), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n444), .A2(new_n446), .A3(new_n247), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n247), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT74), .B(new_n442), .C1(new_n447), .C2(new_n448), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT30), .B(new_n442), .C1(new_n447), .C2(new_n448), .ZN(new_n455));
  INV_X1    g254(.A(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(new_n446), .A3(new_n247), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT35), .B1(new_n399), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n277), .B1(new_n274), .B2(new_n272), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n286), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n468), .A2(new_n280), .B1(new_n397), .B2(new_n392), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n454), .A2(new_n472), .A3(new_n460), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n454), .B2(new_n460), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n438), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT90), .B1(new_n433), .B2(new_n434), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n478), .B(new_n427), .C1(new_n415), .C2(new_n423), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n428), .A2(new_n429), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n471), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n454), .A2(new_n472), .A3(new_n460), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n435), .A2(new_n478), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n431), .A2(KEYINPUT90), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n438), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(KEYINPUT91), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n469), .A2(new_n470), .A3(new_n483), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n463), .A3(new_n280), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n392), .A2(new_n397), .A3(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n398), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT79), .B1(new_n412), .B2(new_n413), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n409), .A2(new_n406), .A3(new_n410), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n421), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT88), .B1(new_n500), .B2(new_n403), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n402), .B1(new_n411), .B2(new_n414), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n404), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT39), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT89), .B1(new_n418), .B2(new_n404), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT39), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n404), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n506), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n427), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n505), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n475), .A2(new_n480), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n451), .A2(new_n453), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n456), .A2(new_n458), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n518), .A2(KEYINPUT37), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(KEYINPUT37), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n457), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT38), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n482), .B(new_n517), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n525), .A3(new_n288), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n464), .A2(new_n492), .B1(new_n497), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(KEYINPUT41), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(KEYINPUT41), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT14), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT14), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G29gat), .B2(G36gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n536), .A2(KEYINPUT94), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(KEYINPUT94), .B2(new_n536), .ZN(new_n538));
  XOR2_X1   g337(.A(G43gat), .B(G50gat), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n540), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n531), .B2(new_n532), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n544), .A2(new_n541), .A3(new_n536), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  INV_X1    g346(.A(G92gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT106), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(KEYINPUT7), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT106), .A3(G85gat), .A4(G92gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n550), .B(new_n552), .C1(KEYINPUT106), .C2(new_n551), .ZN(new_n553));
  XOR2_X1   g352(.A(G99gat), .B(G106gat), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT107), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n547), .B2(new_n548), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n554), .A2(KEYINPUT107), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n530), .B1(new_n546), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n546), .B2(KEYINPUT95), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n565), .B(KEYINPUT17), .C1(new_n542), .C2(new_n545), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n560), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n316), .B(new_n562), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n564), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(G190gat), .B1(new_n570), .B2(new_n561), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(G218gat), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT105), .ZN(new_n573));
  AOI21_X1  g372(.A(G218gat), .B1(new_n569), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n529), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(new_n529), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(KEYINPUT105), .A3(new_n577), .A4(new_n572), .ZN(new_n578));
  XOR2_X1   g377(.A(G134gat), .B(G162gat), .Z(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n575), .B2(new_n578), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(KEYINPUT100), .ZN(new_n591));
  INV_X1    g390(.A(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G64gat), .ZN(new_n593));
  INV_X1    g392(.A(G64gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G57gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n591), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT101), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT102), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G15gat), .B(G22gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT96), .ZN(new_n615));
  INV_X1    g414(.A(G1gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(KEYINPUT16), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G8gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n598), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(KEYINPUT21), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n611), .A3(new_n606), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n623), .B1(new_n613), .B2(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n585), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n584), .A3(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n583), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n598), .A2(new_n560), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT108), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n568), .A2(new_n597), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n634), .A3(KEYINPUT108), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT10), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n568), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n633), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n635), .A2(new_n637), .ZN(new_n642));
  INV_X1    g441(.A(new_n633), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n644), .A3(new_n648), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT109), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT109), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G169gat), .B(G197gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT93), .ZN(new_n658));
  XOR2_X1   g457(.A(G113gat), .B(G141gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n620), .B1(new_n564), .B2(new_n566), .ZN(new_n664));
  INV_X1    g463(.A(G8gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n619), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n546), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(KEYINPUT18), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n666), .B2(new_n546), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n666), .B2(new_n546), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n669), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n620), .B(new_n671), .C1(new_n545), .C2(new_n542), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT18), .B1(new_n668), .B2(new_n669), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n663), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  INV_X1    g481(.A(new_n663), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n678), .A4(new_n670), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT99), .B(new_n663), .C1(new_n679), .C2(new_n680), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR4_X1    g487(.A1(new_n527), .A2(new_n632), .A3(new_n656), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n439), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n616), .ZN(G1324gat));
  XOR2_X1   g490(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n692));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n486), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT111), .Z(new_n696));
  OAI21_X1  g495(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(KEYINPUT42), .A3(new_n695), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n697), .B(new_n698), .C1(new_n665), .C2(new_n693), .ZN(G1325gat));
  AND3_X1   g498(.A1(new_n392), .A2(new_n397), .A3(KEYINPUT36), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT36), .B1(new_n392), .B2(new_n397), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n689), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n398), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n689), .B2(new_n705), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n689), .A2(new_n288), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT43), .B(G22gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  NOR2_X1   g508(.A1(new_n527), .A2(new_n583), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n631), .A2(new_n656), .A3(new_n688), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n439), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n531), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n526), .A2(new_n702), .A3(new_n493), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n483), .A2(new_n470), .A3(new_n491), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n399), .ZN(new_n718));
  INV_X1    g517(.A(new_n463), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n470), .B1(new_n469), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT112), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n464), .A2(new_n492), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(new_n716), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n583), .A2(KEYINPUT44), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n527), .B2(new_n583), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n711), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n439), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n532), .A3(new_n475), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n486), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n730), .A2(new_n737), .A3(new_n702), .ZN(new_n738));
  AOI21_X1  g537(.A(G43gat), .B1(new_n712), .B2(new_n398), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g540(.A(new_n712), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(G50gat), .A3(new_n288), .ZN(new_n743));
  INV_X1    g542(.A(new_n288), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n744), .A3(new_n711), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(G50gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n722), .A2(new_n725), .ZN(new_n748));
  INV_X1    g547(.A(new_n688), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n748), .A2(new_n632), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n656), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n439), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n592), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n751), .A2(new_n486), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  OAI21_X1  g557(.A(G71gat), .B1(new_n751), .B2(new_n702), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n704), .A2(new_n655), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n750), .A2(new_n586), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g562(.A1(new_n751), .A2(new_n288), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n587), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n527), .B2(new_n583), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n575), .A2(new_n578), .ZN(new_n772));
  INV_X1    g571(.A(new_n579), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n580), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n721), .A2(KEYINPUT113), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n628), .A2(new_n630), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n688), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n769), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n768), .B(new_n781), .C1(new_n771), .C2(new_n776), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n547), .A3(new_n713), .A4(new_n656), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n778), .A2(new_n656), .A3(new_n688), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n727), .B2(new_n728), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n439), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(G1336gat));
  NOR3_X1   g590(.A1(new_n655), .A2(G92gat), .A3(new_n486), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT115), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n548), .B1(new_n788), .B2(new_n475), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n794), .A2(KEYINPUT52), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n785), .A2(new_n799), .A3(new_n760), .ZN(new_n800));
  OAI21_X1  g599(.A(G99gat), .B1(new_n789), .B2(new_n702), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1338gat));
  AOI211_X1 g601(.A(new_n770), .B(new_n583), .C1(new_n723), .C2(new_n716), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(new_n721), .B2(new_n775), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n782), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n768), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n777), .A2(new_n769), .A3(new_n782), .ZN(new_n807));
  INV_X1    g606(.A(G106gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n744), .A2(new_n656), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT117), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n788), .A2(new_n744), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n815), .B2(G106gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT118), .A4(new_n814), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n783), .A2(new_n784), .A3(new_n809), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n808), .B1(new_n788), .B2(new_n744), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT53), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(KEYINPUT53), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n828), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n673), .A2(new_n677), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n675), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n668), .A2(new_n669), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n662), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n679), .A2(new_n680), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n683), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n654), .A3(new_n652), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n643), .B(new_n639), .C1(new_n642), .C2(KEYINPUT10), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n641), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n633), .C1(new_n638), .C2(new_n640), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n649), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n641), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n651), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n836), .B1(new_n847), .B2(new_n688), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n583), .ZN(new_n849));
  INV_X1    g648(.A(new_n847), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n775), .A2(new_n835), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n631), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n583), .A2(new_n631), .A3(new_n655), .A4(new_n688), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n439), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n399), .A2(new_n475), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n749), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n855), .A2(new_n744), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n475), .A2(new_n439), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n704), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n688), .A2(new_n342), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n859), .B2(new_n656), .ZN(new_n867));
  INV_X1    g666(.A(new_n863), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n704), .A2(new_n655), .A3(new_n340), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n859), .A2(new_n348), .A3(new_n631), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n863), .A2(new_n704), .A3(new_n778), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n348), .ZN(G1342gat));
  NOR3_X1   g672(.A1(new_n858), .A2(G134gat), .A3(new_n583), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT56), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n863), .A2(new_n704), .A3(new_n583), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n346), .B2(new_n876), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n700), .A2(new_n288), .A3(new_n701), .A4(new_n475), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n208), .B1(new_n879), .B2(new_n688), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n835), .A2(new_n843), .A3(new_n651), .A4(new_n846), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n580), .B2(new_n774), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n583), .B2(new_n848), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n853), .B1(new_n883), .B2(new_n631), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n744), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n702), .A2(new_n862), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n846), .A2(new_n651), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT55), .B1(new_n844), .B2(new_n845), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n843), .A2(KEYINPUT119), .A3(new_n651), .A4(new_n846), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n749), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n775), .B1(new_n893), .B2(new_n836), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n778), .B1(new_n894), .B2(new_n882), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n854), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n288), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n886), .B(new_n887), .C1(new_n899), .C2(new_n885), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n688), .A2(new_n208), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n880), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(new_n879), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n205), .A3(new_n656), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n884), .A2(new_n909), .A3(KEYINPUT57), .A4(new_n744), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT57), .B(new_n744), .C1(new_n852), .C2(new_n854), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n288), .B1(new_n895), .B2(new_n853), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n910), .B(new_n912), .C1(new_n913), .C2(KEYINPUT57), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n656), .A3(new_n887), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n205), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n656), .A4(new_n887), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n908), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n908), .A2(G148gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n900), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n656), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n907), .B1(new_n919), .B2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n906), .B2(new_n631), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n631), .A2(G155gat), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT123), .Z(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n921), .B2(new_n926), .ZN(G1346gat));
  AOI21_X1  g726(.A(G162gat), .B1(new_n906), .B2(new_n775), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n775), .A2(G162gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n921), .B2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n713), .A2(new_n486), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n861), .A2(new_n398), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n688), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n884), .A2(new_n439), .A3(new_n469), .A4(new_n475), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n688), .A2(G169gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  NOR3_X1   g739(.A1(new_n932), .A2(new_n292), .A3(new_n655), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n935), .A2(new_n656), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n292), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n932), .B2(new_n778), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n631), .A2(new_n328), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n934), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n932), .B2(new_n583), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n935), .A2(new_n327), .A3(new_n775), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1351gat));
  NAND3_X1  g750(.A1(new_n702), .A2(new_n744), .A3(new_n475), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT126), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n855), .A2(new_n713), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n749), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n702), .A2(new_n931), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n914), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n749), .A2(G197gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  NOR2_X1   g760(.A1(new_n655), .A2(G204gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  NAND3_X1  g763(.A1(new_n914), .A2(new_n656), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n966), .A3(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n237), .A3(new_n631), .ZN(new_n972));
  OAI21_X1  g771(.A(G211gat), .B1(new_n958), .B2(new_n778), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n958), .B2(new_n583), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n954), .A2(new_n238), .A3(new_n775), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


