

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n524), .B(KEYINPUT17), .ZN(n526) );
  XNOR2_X2 U555 ( .A(n526), .B(n525), .ZN(n607) );
  NOR2_X1 U556 ( .A1(n793), .A2(n776), .ZN(n520) );
  INV_X1 U557 ( .A(n892), .ZN(n776) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n793), .ZN(n768) );
  AND2_X1 U559 ( .A1(n777), .A2(n520), .ZN(n778) );
  INV_X1 U560 ( .A(n708), .ZN(n710) );
  INV_X1 U561 ( .A(KEYINPUT66), .ZN(n524) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n638) );
  NOR2_X1 U565 ( .A1(n627), .A2(G651), .ZN(n645) );
  XNOR2_X1 U566 ( .A(n529), .B(KEYINPUT86), .ZN(n533) );
  INV_X1 U567 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n521), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n522), .B(KEYINPUT65), .ZN(n675) );
  NAND2_X1 U570 ( .A1(n675), .A2(G102), .ZN(n523) );
  XOR2_X1 U571 ( .A(n523), .B(KEYINPUT85), .Z(n528) );
  NAND2_X1 U572 ( .A1(G138), .A2(n607), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n521), .A2(G2104), .ZN(n978) );
  NAND2_X1 U575 ( .A1(G126), .A2(n978), .ZN(n531) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n979) );
  NAND2_X1 U577 ( .A1(G114), .A2(n979), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U579 ( .A1(n533), .A2(n532), .ZN(G164) );
  AND2_X1 U580 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U581 ( .A(G57), .ZN(G237) );
  INV_X1 U582 ( .A(G69), .ZN(G235) );
  INV_X1 U583 ( .A(G108), .ZN(G238) );
  INV_X1 U584 ( .A(G120), .ZN(G236) );
  INV_X1 U585 ( .A(G82), .ZN(G220) );
  NAND2_X1 U586 ( .A1(G88), .A2(n638), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  INV_X1 U588 ( .A(G651), .ZN(n536) );
  NOR2_X1 U589 ( .A1(n627), .A2(n536), .ZN(n641) );
  NAND2_X1 U590 ( .A1(G75), .A2(n641), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G543), .A2(n536), .ZN(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n537) );
  XNOR2_X1 U594 ( .A(n538), .B(n537), .ZN(n637) );
  NAND2_X1 U595 ( .A1(G62), .A2(n637), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G50), .A2(n645), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U598 ( .A1(n542), .A2(n541), .ZN(G166) );
  NAND2_X1 U599 ( .A1(n645), .A2(G51), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT77), .B(n543), .Z(n545) );
  NAND2_X1 U601 ( .A1(n637), .A2(G63), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(KEYINPUT6), .B(n546), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G89), .A2(n638), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT4), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT76), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G76), .A2(n641), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(n551), .B(KEYINPUT5), .Z(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT78), .B(n554), .Z(n555) );
  XNOR2_X1 U612 ( .A(KEYINPUT7), .B(n555), .ZN(G168) );
  XOR2_X1 U613 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n556) );
  XOR2_X1 U615 ( .A(n556), .B(KEYINPUT10), .Z(n1029) );
  NAND2_X1 U616 ( .A1(n1029), .A2(G567), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U618 ( .A1(n645), .A2(G43), .ZN(n558) );
  XNOR2_X1 U619 ( .A(KEYINPUT74), .B(n558), .ZN(n568) );
  XNOR2_X1 U620 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n638), .A2(G81), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G68), .A2(n641), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n637), .A2(G56), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n1008) );
  INV_X1 U630 ( .A(G860), .ZN(n598) );
  OR2_X1 U631 ( .A1(n1008), .A2(n598), .ZN(G153) );
  NAND2_X1 U632 ( .A1(G90), .A2(n638), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G77), .A2(n641), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT9), .B(n571), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G64), .A2(n637), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G52), .A2(n645), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT69), .B(n574), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(G301) );
  INV_X1 U641 ( .A(G301), .ZN(G171) );
  NAND2_X1 U642 ( .A1(G868), .A2(G171), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G66), .A2(n637), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G92), .A2(n638), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G79), .A2(n641), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G54), .A2(n645), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(KEYINPUT15), .B(n583), .ZN(n726) );
  INV_X1 U651 ( .A(n726), .ZN(n1005) );
  INV_X1 U652 ( .A(G868), .ZN(n657) );
  NAND2_X1 U653 ( .A1(n1005), .A2(n657), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U656 ( .A1(n645), .A2(G53), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT70), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G65), .A2(n637), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n590), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G91), .A2(n638), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G78), .A2(n641), .ZN(n591) );
  AND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n657), .ZN(n595) );
  XOR2_X1 U666 ( .A(KEYINPUT79), .B(n595), .Z(n597) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n1005), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n1008), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G868), .A2(n1005), .ZN(n601) );
  NOR2_X1 U674 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n978), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  BUF_X1 U678 ( .A(n675), .Z(n982) );
  NAND2_X1 U679 ( .A1(n982), .A2(G99), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n979), .A2(G111), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G135), .A2(n607), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n991) );
  XNOR2_X1 U685 ( .A(G2096), .B(n991), .ZN(n612) );
  INV_X1 U686 ( .A(G2100), .ZN(n961) );
  NAND2_X1 U687 ( .A1(n612), .A2(n961), .ZN(G156) );
  NAND2_X1 U688 ( .A1(G93), .A2(n638), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT80), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n637), .A2(G67), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT82), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G55), .A2(n645), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G80), .A2(n641), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n656) );
  NAND2_X1 U698 ( .A1(G559), .A2(n1005), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(n1008), .ZN(n654) );
  NOR2_X1 U700 ( .A1(G860), .A2(n654), .ZN(n623) );
  XOR2_X1 U701 ( .A(n656), .B(n623), .Z(G145) );
  NAND2_X1 U702 ( .A1(G49), .A2(n645), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n637), .A2(n626), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U708 ( .A1(n638), .A2(G85), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n637), .A2(G60), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G72), .A2(n641), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G47), .A2(n645), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U715 ( .A(KEYINPUT68), .B(n636), .Z(G290) );
  NAND2_X1 U716 ( .A1(G61), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G86), .A2(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n645), .A2(G48), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(G305) );
  XOR2_X1 U724 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n648) );
  XNOR2_X1 U725 ( .A(n656), .B(n648), .ZN(n649) );
  XNOR2_X1 U726 ( .A(G288), .B(n649), .ZN(n651) );
  XOR2_X1 U727 ( .A(G290), .B(G299), .Z(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U729 ( .A(n652), .B(G166), .Z(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G305), .ZN(n1004) );
  XNOR2_X1 U731 ( .A(n654), .B(n1004), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n655), .A2(G868), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U741 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U742 ( .A1(G219), .A2(G220), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U744 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G96), .A2(n666), .ZN(n953) );
  NAND2_X1 U746 ( .A1(n953), .A2(G2106), .ZN(n671) );
  NOR2_X1 U747 ( .A1(G236), .A2(G238), .ZN(n668) );
  NOR2_X1 U748 ( .A1(G235), .A2(G237), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U750 ( .A(KEYINPUT84), .B(n669), .ZN(n954) );
  NAND2_X1 U751 ( .A1(n954), .A2(G567), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(n955) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n955), .A2(n672), .ZN(n822) );
  NAND2_X1 U755 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(n979), .A2(G113), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G137), .A2(n607), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n674), .A2(n673), .ZN(n680) );
  NAND2_X1 U759 ( .A1(G101), .A2(n675), .ZN(n676) );
  XOR2_X1 U760 ( .A(KEYINPUT23), .B(n676), .Z(n678) );
  NAND2_X1 U761 ( .A1(n978), .A2(G125), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U763 ( .A1(n680), .A2(n679), .ZN(G160) );
  INV_X1 U764 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U765 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n818) );
  XNOR2_X1 U766 ( .A(G1986), .B(G290), .ZN(n884) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n708), .A2(n709), .ZN(n681) );
  XOR2_X1 U769 ( .A(KEYINPUT87), .B(n681), .Z(n813) );
  NAND2_X1 U770 ( .A1(n884), .A2(n813), .ZN(n800) );
  NAND2_X1 U771 ( .A1(G104), .A2(n982), .ZN(n683) );
  NAND2_X1 U772 ( .A1(G140), .A2(n607), .ZN(n682) );
  NAND2_X1 U773 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n684), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G128), .A2(n978), .ZN(n686) );
  NAND2_X1 U776 ( .A1(G116), .A2(n979), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U778 ( .A(KEYINPUT88), .B(n687), .Z(n688) );
  XNOR2_X1 U779 ( .A(KEYINPUT35), .B(n688), .ZN(n689) );
  NOR2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U781 ( .A(KEYINPUT36), .B(n691), .Z(n992) );
  XOR2_X1 U782 ( .A(G2067), .B(KEYINPUT37), .Z(n810) );
  AND2_X1 U783 ( .A1(n992), .A2(n810), .ZN(n944) );
  NAND2_X1 U784 ( .A1(n813), .A2(n944), .ZN(n808) );
  NAND2_X1 U785 ( .A1(n979), .A2(G117), .ZN(n693) );
  NAND2_X1 U786 ( .A1(G141), .A2(n607), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G105), .A2(n982), .ZN(n694) );
  XNOR2_X1 U789 ( .A(n694), .B(KEYINPUT38), .ZN(n695) );
  XNOR2_X1 U790 ( .A(n695), .B(KEYINPUT89), .ZN(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n978), .A2(G129), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n988) );
  AND2_X1 U794 ( .A1(n988), .A2(G1996), .ZN(n935) );
  NAND2_X1 U795 ( .A1(n978), .A2(G119), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G131), .A2(n607), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U798 ( .A1(G95), .A2(n982), .ZN(n703) );
  NAND2_X1 U799 ( .A1(G107), .A2(n979), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n997) );
  INV_X1 U802 ( .A(G1991), .ZN(n853) );
  NOR2_X1 U803 ( .A1(n997), .A2(n853), .ZN(n933) );
  OR2_X1 U804 ( .A1(n935), .A2(n933), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n706), .A2(n813), .ZN(n801) );
  NAND2_X1 U806 ( .A1(n808), .A2(n801), .ZN(n707) );
  XNOR2_X1 U807 ( .A(KEYINPUT90), .B(n707), .ZN(n798) );
  NOR2_X2 U808 ( .A1(n710), .A2(n709), .ZN(n741) );
  NAND2_X1 U809 ( .A1(G2072), .A2(n741), .ZN(n711) );
  XNOR2_X1 U810 ( .A(n711), .B(KEYINPUT27), .ZN(n712) );
  XNOR2_X1 U811 ( .A(n712), .B(KEYINPUT94), .ZN(n714) );
  INV_X1 U812 ( .A(G1956), .ZN(n887) );
  NOR2_X1 U813 ( .A1(n741), .A2(n887), .ZN(n713) );
  NOR2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n717) );
  INV_X1 U815 ( .A(G299), .ZN(n716) );
  OR2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n715) );
  XNOR2_X1 U817 ( .A(n715), .B(KEYINPUT28), .ZN(n734) );
  NAND2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n732) );
  NOR2_X1 U819 ( .A1(n741), .A2(G1348), .ZN(n719) );
  INV_X1 U820 ( .A(n741), .ZN(n757) );
  NOR2_X1 U821 ( .A1(G2067), .A2(n757), .ZN(n718) );
  NOR2_X1 U822 ( .A1(n719), .A2(n718), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n726), .A2(n727), .ZN(n725) );
  AND2_X1 U824 ( .A1(n741), .A2(G1996), .ZN(n720) );
  XOR2_X1 U825 ( .A(KEYINPUT26), .B(n720), .Z(n723) );
  AND2_X1 U826 ( .A1(n757), .A2(G1341), .ZN(n721) );
  NOR2_X1 U827 ( .A1(n721), .A2(n1008), .ZN(n722) );
  AND2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n729) );
  OR2_X1 U830 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U831 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U832 ( .A(KEYINPUT95), .B(n730), .ZN(n731) );
  NAND2_X1 U833 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n736) );
  XOR2_X1 U835 ( .A(KEYINPUT96), .B(KEYINPUT29), .Z(n735) );
  XNOR2_X1 U836 ( .A(n736), .B(n735), .ZN(n740) );
  INV_X1 U837 ( .A(G1961), .ZN(n969) );
  NAND2_X1 U838 ( .A1(n757), .A2(n969), .ZN(n738) );
  XNOR2_X1 U839 ( .A(G2078), .B(KEYINPUT25), .ZN(n854) );
  NAND2_X1 U840 ( .A1(n741), .A2(n854), .ZN(n737) );
  NAND2_X1 U841 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n749), .A2(G171), .ZN(n739) );
  NAND2_X1 U843 ( .A1(n740), .A2(n739), .ZN(n755) );
  XNOR2_X1 U844 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n753) );
  INV_X1 U845 ( .A(G2084), .ZN(n742) );
  AND2_X1 U846 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U847 ( .A(n743), .B(KEYINPUT92), .ZN(n769) );
  INV_X1 U848 ( .A(n769), .ZN(n744) );
  NAND2_X1 U849 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U850 ( .A1(G8), .A2(n757), .ZN(n793) );
  NOR2_X1 U851 ( .A1(n745), .A2(n768), .ZN(n747) );
  XNOR2_X1 U852 ( .A(KEYINPUT30), .B(KEYINPUT97), .ZN(n746) );
  XNOR2_X1 U853 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U854 ( .A1(n748), .A2(G168), .ZN(n751) );
  NOR2_X1 U855 ( .A1(G171), .A2(n749), .ZN(n750) );
  NOR2_X1 U856 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U857 ( .A(n753), .B(n752), .Z(n754) );
  NAND2_X1 U858 ( .A1(n755), .A2(n754), .ZN(n766) );
  AND2_X1 U859 ( .A1(G286), .A2(G8), .ZN(n756) );
  NAND2_X1 U860 ( .A1(n766), .A2(n756), .ZN(n764) );
  INV_X1 U861 ( .A(G8), .ZN(n762) );
  NOR2_X1 U862 ( .A1(G1971), .A2(n793), .ZN(n759) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U864 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U865 ( .A1(n760), .A2(G303), .ZN(n761) );
  OR2_X1 U866 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U867 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U868 ( .A(n765), .B(KEYINPUT32), .ZN(n774) );
  INV_X1 U869 ( .A(n766), .ZN(n767) );
  NOR2_X1 U870 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U871 ( .A1(G8), .A2(n769), .ZN(n770) );
  XOR2_X1 U872 ( .A(KEYINPUT93), .B(n770), .Z(n771) );
  NAND2_X1 U873 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U874 ( .A1(n774), .A2(n773), .ZN(n786) );
  NOR2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n894) );
  NOR2_X1 U876 ( .A1(G1971), .A2(G303), .ZN(n890) );
  NOR2_X1 U877 ( .A1(n894), .A2(n890), .ZN(n775) );
  NAND2_X1 U878 ( .A1(n786), .A2(n775), .ZN(n777) );
  NAND2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n892) );
  XNOR2_X1 U880 ( .A(n778), .B(KEYINPUT64), .ZN(n779) );
  NOR2_X1 U881 ( .A1(KEYINPUT33), .A2(n779), .ZN(n782) );
  NAND2_X1 U882 ( .A1(n894), .A2(KEYINPUT33), .ZN(n780) );
  NOR2_X1 U883 ( .A1(n780), .A2(n793), .ZN(n781) );
  NOR2_X1 U884 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U885 ( .A(G1981), .B(G305), .Z(n880) );
  NAND2_X1 U886 ( .A1(n783), .A2(n880), .ZN(n790) );
  NAND2_X1 U887 ( .A1(G8), .A2(G166), .ZN(n784) );
  NOR2_X1 U888 ( .A1(G2090), .A2(n784), .ZN(n785) );
  XNOR2_X1 U889 ( .A(n785), .B(KEYINPUT99), .ZN(n787) );
  NAND2_X1 U890 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U891 ( .A1(n788), .A2(n793), .ZN(n789) );
  NAND2_X1 U892 ( .A1(n790), .A2(n789), .ZN(n796) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XNOR2_X1 U894 ( .A(n791), .B(KEYINPUT24), .ZN(n792) );
  XNOR2_X1 U895 ( .A(n792), .B(KEYINPUT91), .ZN(n794) );
  NOR2_X1 U896 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U897 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n816) );
  INV_X1 U900 ( .A(n801), .ZN(n804) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n802) );
  AND2_X1 U902 ( .A1(n853), .A2(n997), .ZN(n934) );
  NOR2_X1 U903 ( .A1(n802), .A2(n934), .ZN(n803) );
  NOR2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n988), .ZN(n927) );
  NOR2_X1 U906 ( .A1(n805), .A2(n927), .ZN(n806) );
  XNOR2_X1 U907 ( .A(n806), .B(KEYINPUT39), .ZN(n807) );
  XNOR2_X1 U908 ( .A(n807), .B(KEYINPUT100), .ZN(n809) );
  NAND2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n810), .A2(n992), .ZN(n811) );
  XNOR2_X1 U911 ( .A(n811), .B(KEYINPUT101), .ZN(n924) );
  NAND2_X1 U912 ( .A1(n812), .A2(n924), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U916 ( .A1(n1029), .A2(G2106), .ZN(n819) );
  XOR2_X1 U917 ( .A(KEYINPUT105), .B(n819), .Z(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U919 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U921 ( .A1(n822), .A2(n821), .ZN(G188) );
  NAND2_X1 U923 ( .A1(G100), .A2(n982), .ZN(n824) );
  NAND2_X1 U924 ( .A1(G112), .A2(n979), .ZN(n823) );
  NAND2_X1 U925 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U926 ( .A(KEYINPUT108), .B(n825), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G124), .A2(n978), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n826), .B(KEYINPUT44), .ZN(n828) );
  NAND2_X1 U929 ( .A1(G136), .A2(n607), .ZN(n827) );
  NAND2_X1 U930 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X1 U931 ( .A1(n830), .A2(n829), .ZN(G162) );
  XOR2_X1 U932 ( .A(G20), .B(G1956), .Z(n834) );
  XNOR2_X1 U933 ( .A(G1341), .B(G19), .ZN(n832) );
  XNOR2_X1 U934 ( .A(G6), .B(G1981), .ZN(n831) );
  NOR2_X1 U935 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U936 ( .A1(n834), .A2(n833), .ZN(n837) );
  XOR2_X1 U937 ( .A(KEYINPUT59), .B(G1348), .Z(n835) );
  XNOR2_X1 U938 ( .A(G4), .B(n835), .ZN(n836) );
  NOR2_X1 U939 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U940 ( .A(KEYINPUT60), .B(n838), .ZN(n849) );
  XOR2_X1 U941 ( .A(G1966), .B(G21), .Z(n840) );
  XOR2_X1 U942 ( .A(G1961), .B(G5), .Z(n839) );
  NAND2_X1 U943 ( .A1(n840), .A2(n839), .ZN(n847) );
  XNOR2_X1 U944 ( .A(G1971), .B(G22), .ZN(n842) );
  XNOR2_X1 U945 ( .A(G23), .B(G1976), .ZN(n841) );
  NOR2_X1 U946 ( .A1(n842), .A2(n841), .ZN(n844) );
  XOR2_X1 U947 ( .A(G1986), .B(G24), .Z(n843) );
  NAND2_X1 U948 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U949 ( .A(KEYINPUT58), .B(n845), .ZN(n846) );
  NOR2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U951 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n850), .B(KEYINPUT125), .ZN(n851) );
  XOR2_X1 U953 ( .A(KEYINPUT61), .B(n851), .Z(n852) );
  NOR2_X1 U954 ( .A1(G16), .A2(n852), .ZN(n910) );
  XOR2_X1 U955 ( .A(n853), .B(G25), .Z(n865) );
  XOR2_X1 U956 ( .A(n854), .B(G27), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1996), .B(G32), .ZN(n855) );
  NOR2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(KEYINPUT118), .B(n857), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2067), .B(G26), .ZN(n859) );
  XNOR2_X1 U961 ( .A(G33), .B(G2072), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U963 ( .A(KEYINPUT117), .B(n860), .ZN(n861) );
  NOR2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT119), .B(n863), .ZN(n864) );
  NOR2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G28), .A2(n866), .ZN(n867) );
  XNOR2_X1 U968 ( .A(KEYINPUT53), .B(n867), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT120), .B(G34), .Z(n869) );
  XNOR2_X1 U970 ( .A(G2084), .B(KEYINPUT54), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n873) );
  XNOR2_X1 U973 ( .A(G35), .B(G2090), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT55), .B(n874), .ZN(n876) );
  INV_X1 U976 ( .A(G29), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n877), .A2(G11), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT121), .ZN(n908) );
  XNOR2_X1 U980 ( .A(KEYINPUT56), .B(G16), .ZN(n906) );
  XNOR2_X1 U981 ( .A(G1966), .B(KEYINPUT122), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(G168), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n882), .B(KEYINPUT57), .ZN(n886) );
  XOR2_X1 U985 ( .A(n969), .B(G301), .Z(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n889) );
  XOR2_X1 U988 ( .A(n887), .B(G299), .Z(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n904) );
  INV_X1 U990 ( .A(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n902) );
  XOR2_X1 U992 ( .A(n1005), .B(G1348), .Z(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(KEYINPUT123), .ZN(n900) );
  XOR2_X1 U994 ( .A(n894), .B(KEYINPUT124), .Z(n896) );
  NAND2_X1 U995 ( .A1(G1971), .A2(G303), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n898) );
  XNOR2_X1 U997 ( .A(G1341), .B(n1008), .ZN(n897) );
  NOR2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n911), .B(KEYINPUT126), .ZN(n951) );
  XNOR2_X1 U1006 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n946) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n982), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n607), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(G127), .A2(n978), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(G115), .A2(n979), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(KEYINPUT47), .B(n916), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT109), .B(n919), .Z(n993) );
  XOR2_X1 U1016 ( .A(G2072), .B(n993), .Z(n921) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(n922), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n923), .B(KEYINPUT114), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n932) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n928), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n942) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n991), .ZN(n937) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G2084), .B(G160), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT111), .B(n938), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(n946), .B(n945), .ZN(n947) );
  NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n947), .ZN(n948) );
  XOR2_X1 U1038 ( .A(KEYINPUT116), .B(n948), .Z(n949) );
  NAND2_X1 U1039 ( .A1(n949), .A2(G29), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1041 ( .A(KEYINPUT62), .B(n952), .Z(G311) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1043 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(G325) );
  INV_X1 U1045 ( .A(G325), .ZN(G261) );
  INV_X1 U1046 ( .A(n955), .ZN(G319) );
  XOR2_X1 U1047 ( .A(G2096), .B(KEYINPUT43), .Z(n957) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G2072), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n957), .B(n956), .ZN(n958) );
  XOR2_X1 U1050 ( .A(n958), .B(KEYINPUT106), .Z(n960) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G2678), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n960), .B(n959), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(KEYINPUT42), .B(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G2084), .B(G2078), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n965), .B(n964), .ZN(G227) );
  XOR2_X1 U1057 ( .A(G1981), .B(G1966), .Z(n968) );
  INV_X1 U1058 ( .A(G1996), .ZN(n966) );
  XOR2_X1 U1059 ( .A(n966), .B(G1986), .Z(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n971) );
  XOR2_X1 U1062 ( .A(n969), .B(G1956), .Z(n970) );
  XNOR2_X1 U1063 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1064 ( .A(n973), .B(n972), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G2474), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n975), .B(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G1976), .B(n976), .ZN(n977) );
  XOR2_X1 U1068 ( .A(n977), .B(G1991), .Z(G229) );
  NAND2_X1 U1069 ( .A1(G130), .A2(n978), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(G118), .A2(n979), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n987) );
  NAND2_X1 U1072 ( .A1(G106), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(G142), .A2(n607), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1075 ( .A(n985), .B(KEYINPUT45), .Z(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n989), .B(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n991), .B(n990), .ZN(n996) );
  XNOR2_X1 U1079 ( .A(n992), .B(G162), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(n994), .B(n993), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(n996), .B(n995), .ZN(n1002) );
  XOR2_X1 U1082 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n999) );
  XNOR2_X1 U1083 ( .A(G160), .B(n997), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(n999), .B(n998), .ZN(n1000) );
  XOR2_X1 U1085 ( .A(G164), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1086 ( .A(n1002), .B(n1001), .ZN(n1003) );
  NOR2_X1 U1087 ( .A1(G37), .A2(n1003), .ZN(G395) );
  XNOR2_X1 U1088 ( .A(G286), .B(n1004), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(G301), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1090 ( .A(n1007), .B(n1006), .ZN(n1010) );
  XOR2_X1 U1091 ( .A(n1008), .B(KEYINPUT110), .Z(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NOR2_X1 U1093 ( .A1(G37), .A2(n1011), .ZN(G397) );
  XNOR2_X1 U1094 ( .A(G1348), .B(G2446), .ZN(n1021) );
  XOR2_X1 U1095 ( .A(G2454), .B(KEYINPUT104), .Z(n1013) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G2430), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1013), .B(n1012), .ZN(n1017) );
  XOR2_X1 U1098 ( .A(G2443), .B(G2451), .Z(n1015) );
  XNOR2_X1 U1099 ( .A(KEYINPUT103), .B(G2427), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1015), .B(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(n1017), .B(n1016), .Z(n1019) );
  XNOR2_X1 U1102 ( .A(G2435), .B(G2438), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(n1019), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(G14), .ZN(n1028) );
  NAND2_X1 U1106 ( .A1(G319), .A2(n1028), .ZN(n1025) );
  NOR2_X1 U1107 ( .A1(G227), .A2(G229), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT49), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  NOR2_X1 U1110 ( .A1(G395), .A2(G397), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(G225) );
  INV_X1 U1112 ( .A(G225), .ZN(G308) );
  INV_X1 U1113 ( .A(n1028), .ZN(G401) );
  INV_X1 U1114 ( .A(n1029), .ZN(G223) );
endmodule

