//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n188), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT30), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n194), .A2(KEYINPUT65), .A3(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT65), .B1(new_n194), .B2(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n194), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n194), .A2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n193), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n201), .A2(new_n205), .B1(G131), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n208), .B2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(KEYINPUT66), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n212), .A3(new_n214), .A4(new_n209), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n191), .B1(new_n211), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n212), .A3(new_n209), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n216), .A2(new_n212), .A3(KEYINPUT67), .A4(new_n209), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(G131), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n193), .A2(new_n204), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT0), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(KEYINPUT0), .B2(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n230), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n192), .B2(G143), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n194), .A2(KEYINPUT65), .A3(G146), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n198), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n228), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n190), .B1(new_n222), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n202), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n205), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n210), .A2(G131), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n218), .A2(new_n219), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n218), .A2(new_n219), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n248), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n243), .B1(new_n221), .B2(new_n227), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n191), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n228), .A2(new_n244), .B1(new_n211), .B2(new_n221), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n246), .A2(new_n255), .B1(new_n190), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n187), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n245), .A2(new_n190), .A3(new_n252), .ZN(new_n265));
  INV_X1    g079(.A(new_n190), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n253), .B2(new_n254), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT28), .B1(new_n256), .B2(new_n190), .ZN(new_n269));
  INV_X1    g083(.A(new_n262), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT28), .ZN(new_n274));
  INV_X1    g088(.A(new_n269), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n274), .A2(KEYINPUT29), .A3(new_n275), .A4(new_n262), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G472), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n226), .A2(G131), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n225), .A2(new_n281), .B1(new_n217), .B2(new_n220), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT30), .B(new_n252), .C1(new_n282), .C2(new_n243), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n283), .B(new_n266), .C1(new_n256), .C2(KEYINPUT30), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n270), .B1(new_n256), .B2(new_n190), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n284), .A2(KEYINPUT31), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT31), .B1(new_n284), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n295), .B(new_n279), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  INV_X1    g110(.A(G217), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(G234), .B2(new_n277), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G125), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(KEYINPUT70), .A3(G125), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT16), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n192), .A2(KEYINPUT71), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n192), .A2(KEYINPUT71), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n307), .A2(new_n315), .A3(G146), .A4(new_n309), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n202), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n322), .A2(new_n321), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT24), .B(G110), .Z(new_n327));
  AOI22_X1  g141(.A1(new_n325), .A2(G110), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n316), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n310), .A2(G146), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT72), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n192), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n325), .A2(G110), .B1(new_n326), .B2(new_n327), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G221), .A3(G234), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT73), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G137), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n329), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n329), .B2(new_n335), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n277), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT25), .B(new_n277), .C1(new_n341), .C2(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n299), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n329), .A2(new_n335), .ZN(new_n348));
  INV_X1    g162(.A(new_n340), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n329), .A2(new_n335), .A3(new_n340), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n298), .A2(G902), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n294), .A2(new_n296), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n361));
  INV_X1    g175(.A(G113), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G119), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n361), .A2(new_n366), .B1(new_n188), .B2(new_n189), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G104), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT75), .B(G107), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G101), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g193(.A(G101), .B1(new_n373), .B2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n367), .A2(new_n372), .A3(KEYINPUT79), .A4(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n373), .A2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n379), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT4), .A3(G101), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n190), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n360), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(KEYINPUT4), .A2(new_n381), .B1(new_n388), .B2(G101), .ZN(new_n395));
  INV_X1    g209(.A(new_n392), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n266), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n397), .A2(new_n359), .A3(new_n384), .A4(new_n385), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT6), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n360), .C1(new_n386), .C2(new_n393), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n197), .A2(new_n200), .B1(new_n229), .B2(new_n203), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n302), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n244), .B2(new_n302), .ZN(new_n404));
  INV_X1    g218(.A(G224), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G953), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n404), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n405), .B2(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n372), .A2(new_n381), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n367), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n359), .B(KEYINPUT8), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n318), .A2(G116), .ZN(new_n414));
  OAI21_X1  g228(.A(G113), .B1(new_n414), .B2(KEYINPUT5), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n361), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n189), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n417), .A2(new_n418), .B1(new_n189), .B2(new_n188), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n412), .B(new_n413), .C1(new_n411), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n409), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n403), .B(new_n421), .C1(new_n244), .C2(new_n302), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n410), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n423), .B2(new_n398), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n408), .A2(new_n424), .A3(new_n426), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n358), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G237), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n336), .A3(G214), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n194), .ZN(new_n433));
  AOI21_X1  g247(.A(G143), .B1(new_n258), .B2(G214), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n194), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n214), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT17), .A3(G131), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n314), .B2(new_n316), .ZN(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(new_n373), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(KEYINPUT18), .A3(G131), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n438), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n305), .A2(new_n306), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n305), .A2(KEYINPUT82), .A3(new_n306), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(G146), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n451), .B1(new_n456), .B2(new_n333), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n444), .A2(new_n447), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(KEYINPUT19), .A3(new_n455), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n332), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n461), .A3(new_n192), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n310), .A2(G146), .B1(new_n435), .B2(new_n439), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n333), .ZN(new_n465));
  INV_X1    g279(.A(new_n451), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n446), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G475), .A2(G902), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT83), .B1(new_n458), .B2(new_n468), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n314), .A2(new_n316), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n467), .B(new_n446), .C1(new_n475), .C2(new_n443), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n446), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n473), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n447), .B1(new_n444), .B2(new_n457), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n476), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n277), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(G475), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n202), .B2(G143), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n194), .A2(KEYINPUT13), .A3(G128), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n202), .A2(G143), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G134), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n202), .A2(G143), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n492), .A3(new_n208), .ZN(new_n497));
  XNOR2_X1  g311(.A(G116), .B(G122), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n370), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n370), .A2(new_n498), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n494), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n370), .B(new_n498), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n494), .A4(new_n497), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n194), .A2(G128), .ZN(new_n506));
  OAI21_X1  g320(.A(G134), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n497), .A2(new_n507), .B1(new_n370), .B2(new_n498), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n363), .A2(KEYINPUT14), .A3(G122), .ZN(new_n509));
  INV_X1    g323(.A(new_n498), .ZN(new_n510));
  OAI211_X1 g324(.A(G107), .B(new_n509), .C1(new_n510), .C2(KEYINPUT14), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n505), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT9), .B(G234), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n514), .A2(new_n297), .A3(G953), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n501), .A2(new_n502), .B1(new_n511), .B2(new_n508), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n277), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT85), .ZN(new_n521));
  INV_X1    g335(.A(G478), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n513), .A2(new_n516), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n505), .A3(new_n515), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n526), .B1(KEYINPUT15), .B2(new_n522), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n336), .A2(G952), .ZN(new_n532));
  NAND2_X1  g346(.A1(G234), .A2(G237), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT21), .B(G898), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(G902), .A3(G953), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n430), .A2(new_n488), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n514), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n205), .B1(new_n229), .B2(new_n247), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n372), .A2(new_n381), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n248), .B1(new_n381), .B2(new_n372), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n411), .A2(new_n402), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n228), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n544), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n372), .A2(new_n381), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT77), .B(new_n546), .C1(new_n554), .C2(new_n248), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n555), .A2(KEYINPUT12), .A3(new_n228), .A4(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n402), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n559), .A2(new_n554), .B1(new_n546), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n391), .A2(new_n392), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT76), .B1(new_n561), .B2(new_n244), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n563), .B(new_n243), .C1(new_n391), .C2(new_n392), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n282), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G140), .ZN(new_n567));
  INV_X1    g381(.A(G227), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT74), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(new_n554), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n546), .A2(new_n558), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n244), .B1(new_n395), .B2(new_n396), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n563), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n244), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n570), .B1(new_n579), .B2(new_n282), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n228), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n572), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G469), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n543), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n566), .A2(new_n571), .B1(new_n580), .B2(new_n582), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT78), .B(G469), .C1(new_n587), .C2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n570), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n582), .B2(new_n565), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n557), .A2(new_n565), .A3(new_n589), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n585), .B(new_n277), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n541), .A2(new_n542), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n356), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(G101), .Z(G3));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n542), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n288), .A2(new_n277), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT86), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n288), .A2(new_n290), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(KEYINPUT86), .A3(G472), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n355), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT87), .Z(new_n607));
  NAND2_X1  g421(.A1(new_n480), .A2(new_n482), .ZN(new_n608));
  INV_X1    g422(.A(new_n473), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n487), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT90), .B(G478), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n521), .A2(new_n528), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT33), .B1(new_n517), .B2(new_n519), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n524), .A2(new_n616), .A3(new_n525), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n522), .A2(G902), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT89), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT89), .ZN(new_n621));
  INV_X1    g435(.A(new_n619), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n621), .B(new_n622), .C1(new_n615), .C2(new_n617), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n614), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n612), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n428), .A2(KEYINPUT88), .A3(new_n429), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n426), .B1(new_n408), .B2(new_n424), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n358), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n625), .A2(new_n630), .A3(new_n539), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n607), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  OR2_X1    g448(.A1(new_n480), .A2(new_n482), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n487), .B1(new_n635), .B2(new_n608), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n531), .ZN(new_n637));
  INV_X1    g451(.A(new_n630), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n538), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n607), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  AOI21_X1  g457(.A(KEYINPUT25), .B1(new_n352), .B2(new_n277), .ZN(new_n644));
  INV_X1    g458(.A(new_n346), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n298), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n349), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n348), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n329), .A2(new_n349), .A3(new_n335), .A4(new_n647), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n353), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT91), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT91), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n649), .A2(new_n653), .A3(new_n353), .A4(new_n650), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n646), .A2(new_n655), .A3(KEYINPUT92), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT92), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n654), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n657), .B1(new_n347), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n604), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n542), .ZN(new_n662));
  OAI21_X1  g476(.A(G469), .B1(new_n587), .B2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n582), .A2(new_n565), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n570), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n580), .A2(new_n557), .ZN(new_n666));
  AOI21_X1  g480(.A(G902), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n663), .A2(new_n543), .B1(new_n667), .B2(new_n585), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n662), .B1(new_n668), .B2(new_n588), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n661), .A2(new_n669), .A3(new_n541), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT93), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  NAND4_X1  g487(.A1(new_n294), .A2(new_n296), .A3(new_n542), .A4(new_n593), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n537), .A2(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n534), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n636), .A2(new_n531), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n630), .A2(new_n660), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n202), .ZN(G30));
  XNOR2_X1  g496(.A(new_n676), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n669), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT40), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n660), .A2(new_n357), .A3(new_n612), .A4(new_n531), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n428), .A2(new_n429), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT38), .Z(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n270), .B1(new_n284), .B2(new_n265), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n265), .A2(new_n267), .A3(new_n270), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT94), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT94), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n696), .B(new_n693), .C1(new_n257), .C2(new_n270), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n277), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n291), .B2(new_n292), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n690), .A2(new_n691), .A3(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n685), .A2(new_n687), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n194), .ZN(G45));
  AND4_X1   g517(.A1(new_n294), .A2(new_n296), .A3(new_n542), .A4(new_n593), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n656), .A2(new_n659), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n638), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n624), .B(new_n676), .C1(new_n487), .C2(new_n483), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  INV_X1    g524(.A(new_n631), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n277), .B1(new_n590), .B2(new_n591), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n542), .A3(new_n592), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n294), .A2(new_n296), .A3(new_n355), .A4(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n639), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n363), .ZN(G18));
  NAND2_X1  g534(.A1(new_n294), .A2(new_n296), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n488), .A2(new_n540), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(KEYINPUT96), .A3(new_n679), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT96), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n679), .A2(new_n723), .A3(new_n714), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n721), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND4_X1   g544(.A1(new_n612), .A2(new_n531), .A3(new_n626), .A4(new_n629), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n598), .A2(G472), .B1(new_n288), .B2(new_n290), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n355), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n731), .A2(new_n734), .A3(new_n538), .A4(new_n714), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NAND3_X1  g550(.A1(new_n713), .A2(new_n542), .A3(new_n592), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n630), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n705), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT97), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n612), .A2(new_n742), .A3(new_n624), .A4(new_n676), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n740), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n408), .A2(new_n424), .A3(new_n426), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n627), .A3(new_n358), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n749), .A3(new_n542), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n294), .A3(new_n296), .A4(new_n355), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n741), .A2(new_n743), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n753), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n293), .A2(new_n355), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(KEYINPUT42), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  INV_X1    g573(.A(new_n356), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n678), .A3(new_n751), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n488), .A2(new_n624), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT100), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  INV_X1    g580(.A(new_n604), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n660), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT101), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT101), .A3(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n572), .A2(new_n583), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n585), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT98), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n776), .B2(new_n775), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(KEYINPUT98), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n782), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n592), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n785), .B2(KEYINPUT99), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT99), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n787), .A3(new_n592), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n662), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n790));
  INV_X1    g604(.A(new_n749), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n774), .A2(new_n789), .A3(new_n683), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(new_n707), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n791), .A2(new_n355), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n721), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n300), .ZN(G42));
  NAND2_X1  g615(.A1(new_n713), .A2(new_n592), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT106), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n662), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n799), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n534), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n766), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n734), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n791), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(KEYINPUT108), .A2(KEYINPUT50), .ZN(new_n813));
  OR4_X1    g627(.A1(new_n357), .A2(new_n690), .A3(new_n737), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT108), .B1(KEYINPUT107), .B2(KEYINPUT50), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n737), .A2(new_n791), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n819), .A2(new_n605), .A3(new_n534), .A4(new_n700), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(new_n612), .A3(new_n624), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n809), .A2(new_n740), .A3(new_n818), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n822), .B2(new_n824), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n817), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n812), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n809), .A2(new_n756), .A3(new_n818), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT48), .Z(new_n832));
  INV_X1    g646(.A(new_n738), .ZN(new_n833));
  OAI221_X1 g647(.A(new_n532), .B1(new_n625), .B2(new_n821), .C1(new_n810), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n824), .A4(new_n822), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n807), .B2(new_n811), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n830), .B(new_n835), .C1(new_n839), .C2(KEYINPUT51), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT103), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n662), .B1(new_n663), .B2(new_n592), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n705), .A3(new_n732), .A4(new_n749), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n753), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n750), .A2(new_n739), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT103), .A3(new_n741), .A4(new_n743), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n531), .B1(new_n534), .B2(new_n675), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n636), .A2(new_n705), .A3(new_n749), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n669), .A2(new_n849), .A3(new_n294), .A4(new_n296), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n758), .A2(new_n761), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n715), .B1(new_n711), .B2(new_n639), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n735), .B1(new_n356), .B2(new_n594), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n430), .A2(new_n538), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n488), .A2(new_n531), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n625), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n541), .A2(new_n542), .A3(new_n593), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n606), .A2(new_n858), .B1(new_n859), .B2(new_n661), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n729), .A2(new_n853), .A3(new_n855), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n706), .A2(new_n677), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n739), .A2(new_n737), .A3(new_n630), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n704), .A2(new_n863), .B1(new_n755), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n646), .A2(new_n655), .A3(new_n676), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n842), .A2(new_n700), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n612), .A2(new_n531), .A3(new_n626), .A4(new_n629), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n704), .B2(new_n708), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n744), .B1(new_n674), .B2(new_n680), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n731), .A2(new_n700), .A3(new_n842), .A4(new_n866), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n679), .A2(new_n795), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n674), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT52), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT104), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT104), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n862), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT105), .B(KEYINPUT53), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n844), .A2(new_n846), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n850), .B1(new_n677), .B2(new_n752), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n852), .B1(new_n728), .B2(new_n725), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n858), .A2(new_n669), .A3(new_n767), .A4(new_n355), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n670), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n854), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n888), .A2(new_n889), .A3(new_n758), .A4(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n878), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n884), .A2(new_n885), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n880), .B1(new_n872), .B2(new_n877), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n883), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n881), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n893), .B2(new_n878), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n885), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n840), .A2(new_n905), .B1(G952), .B2(G953), .ZN(new_n906));
  OR4_X1    g720(.A1(new_n605), .A2(new_n763), .A3(new_n662), .A4(new_n358), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT102), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n690), .A2(new_n700), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n802), .B(KEYINPUT49), .Z(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(G75));
  OR3_X1    g728(.A1(new_n336), .A2(KEYINPUT114), .A3(G952), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT114), .B1(new_n336), .B2(G952), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT115), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n901), .B1(new_n900), .B2(new_n881), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n895), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n277), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n399), .A2(new_n401), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n407), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n919), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(KEYINPUT112), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT112), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n921), .B2(new_n277), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n427), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT113), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n928), .B1(new_n933), .B2(new_n935), .ZN(G51));
  AND2_X1   g750(.A1(new_n929), .A2(new_n931), .ZN(new_n937));
  INV_X1    g751(.A(new_n781), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT54), .B1(new_n920), .B2(new_n895), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n941), .A3(new_n897), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n884), .A2(new_n896), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n782), .B(KEYINPUT57), .Z(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n590), .B2(new_n591), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n917), .B1(new_n939), .B2(new_n947), .ZN(G54));
  NAND2_X1  g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT117), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n937), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n474), .A3(new_n479), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n474), .A2(new_n479), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n937), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n917), .B1(new_n952), .B2(new_n954), .ZN(G60));
  INV_X1    g769(.A(new_n618), .ZN(new_n956));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n942), .A2(new_n944), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT118), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n942), .A2(KEYINPUT118), .A3(new_n944), .A4(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n958), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n898), .B2(new_n904), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n918), .B1(new_n966), .B2(new_n956), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT119), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT119), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n964), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT121), .ZN(new_n974));
  XOR2_X1   g788(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n943), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n352), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n918), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT61), .B1(new_n979), .B2(KEYINPUT122), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n649), .A2(new_n650), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(new_n977), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G66));
  AOI21_X1  g797(.A(new_n336), .B1(new_n536), .B2(G224), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n861), .B2(new_n336), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n924), .B1(G898), .B2(new_n336), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(G69));
  INV_X1    g801(.A(G900), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n568), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n255), .A2(new_n283), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT123), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n459), .A2(new_n461), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n756), .A2(new_n731), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n774), .B2(new_n792), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n789), .A2(new_n683), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n709), .A2(new_n758), .A3(new_n761), .A4(new_n865), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n336), .B1(new_n1000), .B2(new_n800), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n988), .A2(G953), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT126), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n994), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n989), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n865), .A2(new_n709), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n702), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n791), .B1(new_n625), .B2(new_n857), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n760), .A2(new_n669), .A3(new_n683), .A4(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1009), .A2(new_n793), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n336), .B1(new_n1012), .B2(new_n800), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n994), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1003), .ZN(new_n1015));
  INV_X1    g829(.A(new_n800), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n998), .A3(new_n999), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n1017), .B2(new_n336), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n1018), .B2(new_n994), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1006), .B(new_n1019), .ZN(G72));
  AND2_X1   g834(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1021));
  INV_X1    g835(.A(new_n861), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1021), .A2(new_n1016), .A3(new_n793), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n692), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1025), .B1(new_n1017), .B2(new_n861), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1030), .A2(new_n270), .A3(new_n257), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n902), .A2(new_n903), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n284), .A2(new_n285), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n257), .A2(new_n262), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1032), .B(new_n1025), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1031), .A2(new_n915), .A3(new_n916), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1029), .A2(new_n1036), .ZN(G57));
endmodule


