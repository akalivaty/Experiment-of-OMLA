//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  OR2_X1    g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n206), .B1(new_n203), .B2(KEYINPUT2), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n215));
  INV_X1    g014(.A(new_n203), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n202), .A2(KEYINPUT74), .A3(new_n203), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n210), .A2(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n208), .A2(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n214), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G211gat), .A2(G218gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n225), .B1(new_n242), .B2(new_n228), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n219), .A2(new_n223), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n204), .A2(new_n215), .B1(KEYINPUT2), .B2(new_n203), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT73), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n223), .A3(new_n207), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n246), .A2(new_n247), .B1(new_n249), .B2(new_n205), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n214), .A2(new_n224), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n237), .B2(new_n241), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n252), .B(new_n253), .C1(new_n225), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n244), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G228gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n214), .A2(new_n224), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n214), .B2(new_n224), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n244), .B(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT80), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n265), .A3(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(G22gat), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n258), .A2(new_n265), .A3(new_n276), .A4(new_n271), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n266), .A2(new_n272), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n275), .A2(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT71), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT68), .B(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  AND2_X1   g088(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n288), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OR3_X1    g099(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n298), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT70), .B1(new_n299), .B2(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT27), .B(G183gat), .Z(new_n305));
  OAI21_X1  g104(.A(KEYINPUT28), .B1(new_n305), .B2(new_n287), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n295), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n299), .B2(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n314), .B(new_n315), .C1(G183gat), .C2(G190gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n297), .B1(KEYINPUT23), .B2(new_n299), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n290), .A2(new_n291), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n287), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n319), .B1(new_n309), .B2(new_n311), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT23), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n296), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT66), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT66), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n332), .A3(new_n296), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n325), .A2(new_n326), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n320), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n320), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n307), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n286), .B1(new_n338), .B2(new_n228), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n334), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n340), .A2(new_n307), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(new_n284), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n243), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT37), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n286), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n284), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n242), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n344), .B1(new_n343), .B2(new_n347), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n283), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n228), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n342), .B1(new_n356), .B2(new_n285), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n355), .B(new_n347), .C1(new_n357), .C2(new_n242), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G1gat), .B(G29gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n261), .B2(new_n262), .ZN(new_n364));
  XNOR2_X1  g163(.A(G127gat), .B(G134gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G113gat), .B(G120gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(KEYINPUT1), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n365), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n364), .A2(new_n373), .A3(new_n227), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n250), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n214), .A2(new_n224), .A3(new_n368), .A4(new_n371), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n373), .B1(new_n261), .B2(new_n262), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n378), .ZN(new_n384));
  INV_X1    g183(.A(new_n375), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n377), .B2(new_n379), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n382), .A3(new_n375), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n363), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n381), .A2(new_n386), .ZN(new_n396));
  INV_X1    g195(.A(new_n363), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n397), .C1(new_n392), .C2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n345), .A2(new_n243), .A3(new_n346), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT37), .B(new_n401), .C1(new_n357), .C2(new_n243), .ZN(new_n402));
  INV_X1    g201(.A(new_n283), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n348), .A2(new_n402), .A3(new_n351), .A4(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT6), .B(new_n363), .C1(new_n387), .C2(new_n394), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n358), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n355), .A4(new_n347), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n307), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n340), .A2(KEYINPUT69), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n320), .A2(new_n334), .A3(new_n335), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n285), .B1(new_n414), .B2(KEYINPUT29), .ZN(new_n415));
  INV_X1    g214(.A(new_n342), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n242), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n347), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n351), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT72), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(new_n351), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n410), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT40), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n380), .A2(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n389), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n374), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n385), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n397), .B1(new_n428), .B2(KEYINPUT39), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n383), .A2(new_n375), .A3(new_n378), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT39), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT81), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n433), .A3(KEYINPUT39), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n375), .B1(new_n426), .B2(new_n374), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n424), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n363), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(KEYINPUT40), .C1(new_n436), .C2(new_n435), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n395), .A3(new_n441), .ZN(new_n442));
  OAI221_X1 g241(.A(new_n282), .B1(new_n359), .B2(new_n406), .C1(new_n423), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n338), .A2(new_n373), .ZN(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT64), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n372), .B(new_n307), .C1(new_n336), .C2(new_n337), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT34), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n444), .B2(new_n448), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(KEYINPUT33), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n444), .A2(new_n448), .ZN(new_n459));
  AOI221_X4 g258(.A(new_n456), .B1(KEYINPUT33), .B2(new_n453), .C1(new_n459), .C2(new_n446), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n450), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n412), .A2(new_n413), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n372), .B1(new_n462), .B2(new_n307), .ZN(new_n463));
  INV_X1    g262(.A(new_n448), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n446), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(new_n453), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n455), .A2(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n449), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(KEYINPUT36), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n458), .A2(new_n450), .A3(new_n460), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n400), .A2(new_n405), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n408), .A2(new_n409), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n420), .A2(new_n422), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n282), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n474), .A2(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n282), .A2(new_n461), .A3(new_n473), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n282), .A2(new_n461), .A3(new_n473), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT35), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n443), .A2(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G113gat), .B(G141gat), .ZN(new_n492));
  INV_X1    g291(.A(G197gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT11), .B(G169gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT12), .ZN(new_n497));
  XOR2_X1   g296(.A(G15gat), .B(G22gat), .Z(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  AOI21_X1  g300(.A(G8gat), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT16), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(G1gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n500), .B1(new_n504), .B2(new_n498), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n502), .B(new_n505), .Z(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G43gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n512), .B2(G50gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n268), .A2(G43gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  OR4_X1    g317(.A1(KEYINPUT85), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n515), .A2(new_n517), .A3(new_n518), .A4(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n528), .A3(new_n520), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(new_n518), .C1(new_n528), .C2(new_n524), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n516), .A4(new_n508), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n506), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT88), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n502), .B(new_n505), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n527), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n534), .A2(new_n535), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n497), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n536), .A2(new_n531), .A3(new_n527), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT13), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n535), .A4(new_n543), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n546), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n548), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  INV_X1    g357(.A(G71gat), .ZN(new_n559));
  INV_X1    g358(.A(G78gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n562));
  XOR2_X1   g361(.A(G57gat), .B(G64gat), .Z(new_n563));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n536), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G183gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT91), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G211gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n577), .B(new_n579), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n576), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT92), .B(G134gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G99gat), .B(G106gat), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT95), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AND2_X1   g388(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  INV_X1    g392(.A(G99gat), .ZN(new_n594));
  INV_X1    g393(.A(G106gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT8), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n592), .B2(new_n596), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n586), .B(new_n588), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n585), .A2(KEYINPUT95), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n596), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT94), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n600), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n606), .A3(new_n586), .A4(new_n588), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n601), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n541), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n532), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n615), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n615), .B2(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n625));
  INV_X1    g424(.A(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n601), .A2(new_n607), .A3(new_n610), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n610), .B1(new_n601), .B2(new_n607), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n632), .A2(new_n541), .B1(new_n532), .B2(new_n608), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n621), .B(new_n620), .C1(new_n633), .C2(new_n618), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n619), .A3(new_n622), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n584), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n627), .B1(new_n623), .B2(new_n624), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n635), .A3(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n583), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n608), .A2(new_n568), .ZN(new_n642));
  INV_X1    g441(.A(new_n568), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n601), .B2(new_n607), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  INV_X1    g449(.A(G233gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n654), .B(new_n660), .C1(new_n645), .C2(new_n653), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n653), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n582), .A2(new_n641), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n491), .A2(new_n557), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n479), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(G8gat), .ZN(new_n672));
  INV_X1    g471(.A(new_n423), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n675), .B2(KEYINPUT42), .ZN(new_n676));
  NOR2_X1   g475(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n503), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  MUX2_X1   g478(.A(new_n672), .B(new_n676), .S(new_n679), .Z(G1325gat));
  NOR2_X1   g479(.A1(new_n476), .A2(new_n477), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n668), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n478), .A2(new_n474), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT101), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n682), .B1(new_n668), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n483), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n582), .A2(new_n665), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n637), .A2(new_n640), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n557), .A3(new_n491), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G29gat), .A3(new_n479), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n691), .A2(new_n556), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n491), .B2(new_n641), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n482), .A2(new_n483), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n282), .B1(new_n423), .B2(new_n442), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n359), .A2(new_n406), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n704), .B(new_n683), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n488), .A2(new_n490), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n692), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n702), .B1(new_n703), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT105), .B(new_n702), .C1(new_n703), .C2(new_n713), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n479), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n719), .ZN(G1328gat));
  OR3_X1    g519(.A1(new_n718), .A2(KEYINPUT106), .A3(new_n423), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT106), .B1(new_n718), .B2(new_n423), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(G36gat), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n698), .A2(G36gat), .A3(new_n423), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT46), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  INV_X1    g526(.A(new_n702), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n692), .B(KEYINPUT104), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n491), .A2(KEYINPUT44), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n710), .B1(new_n709), .B2(new_n692), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n715), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n683), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n727), .B1(new_n735), .B2(new_n512), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n696), .A2(new_n512), .A3(new_n681), .A4(new_n697), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n684), .B1(new_n716), .B2(new_n717), .ZN(new_n738));
  INV_X1    g537(.A(new_n512), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n732), .B2(new_n683), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n737), .A3(KEYINPUT47), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1330gat));
  AOI21_X1  g545(.A(new_n282), .B1(new_n733), .B2(new_n734), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n747), .B2(new_n268), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n282), .B1(new_n698), .B2(KEYINPUT110), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n696), .A2(new_n750), .A3(new_n697), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n268), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n483), .B1(new_n716), .B2(new_n717), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(G50gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G50gat), .B1(new_n732), .B2(new_n282), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n752), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n491), .A2(new_n556), .ZN(new_n762));
  INV_X1    g561(.A(new_n582), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n763), .A2(new_n692), .A3(new_n666), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n669), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n423), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  AOI21_X1  g572(.A(G71gat), .B1(new_n766), .B2(new_n681), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n765), .A2(new_n559), .A3(new_n683), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n765), .A2(new_n282), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT112), .B(G78gat), .Z(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n590), .A2(new_n591), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n582), .A2(new_n556), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n709), .A2(new_n692), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(new_n665), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n782), .B1(new_n787), .B2(new_n669), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n665), .B(new_n783), .C1(new_n730), .C2(new_n731), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n479), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n782), .B2(new_n790), .ZN(G1336gat));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n589), .A3(new_n673), .ZN(new_n792));
  OAI21_X1  g591(.A(G92gat), .B1(new_n789), .B2(new_n423), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n787), .A2(new_n594), .A3(new_n681), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n789), .A2(new_n683), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT113), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n594), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n483), .A2(new_n665), .A3(new_n595), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT114), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  OAI21_X1  g602(.A(G106gat), .B1(new_n789), .B2(new_n282), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  INV_X1    g606(.A(new_n800), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT53), .B1(new_n786), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n804), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1339gat));
  NAND4_X1  g610(.A1(new_n546), .A2(new_n553), .A3(new_n497), .A4(new_n554), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n534), .A2(new_n549), .A3(new_n551), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n535), .B1(new_n534), .B2(new_n543), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n496), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n665), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n660), .B1(new_n662), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n661), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(KEYINPUT116), .A3(new_n825), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n819), .B1(new_n832), .B2(new_n557), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n729), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n830), .A2(new_n828), .A3(new_n831), .A4(new_n818), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n712), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n582), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n667), .A2(new_n556), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g638(.A1(new_n669), .A2(new_n839), .A3(new_n423), .A4(new_n486), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n556), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n665), .ZN(new_n843));
  INV_X1    g642(.A(G120gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n843), .B2(new_n845), .ZN(G1341gat));
  NAND2_X1  g647(.A1(new_n840), .A2(new_n582), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n840), .A2(new_n692), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT56), .B1(new_n851), .B2(G134gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(G134gat), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  INV_X1    g653(.A(G134gat), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n854), .A3(new_n855), .A4(new_n692), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(G1343gat));
  NOR3_X1   g656(.A1(new_n684), .A2(new_n479), .A3(new_n673), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n821), .B(new_n823), .C1(KEYINPUT118), .C2(KEYINPUT55), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n548), .A2(new_n555), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n548), .A2(new_n555), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n661), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n821), .C2(new_n823), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n819), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n641), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n582), .B1(new_n866), .B2(new_n836), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n483), .B1(new_n867), .B2(new_n838), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n859), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n483), .C1(new_n837), .C2(new_n838), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n869), .A2(G141gat), .A3(new_n556), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n483), .B(new_n858), .C1(new_n837), .C2(new_n838), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n208), .B1(new_n873), .B2(new_n557), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT119), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1344gat));
  OAI21_X1  g676(.A(new_n210), .B1(new_n873), .B2(new_n666), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n483), .A2(new_n870), .ZN(new_n879));
  INV_X1    g678(.A(new_n864), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n556), .A2(new_n880), .A3(new_n661), .A4(new_n860), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n692), .B1(new_n881), .B2(new_n819), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n832), .A2(new_n641), .A3(new_n817), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n763), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n838), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n483), .B1(new_n837), .B2(new_n838), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n665), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n858), .A2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n878), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g690(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n892));
  AND2_X1   g691(.A1(new_n869), .A2(new_n871), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n665), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n210), .A2(KEYINPUT59), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n891), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  INV_X1    g695(.A(new_n873), .ZN(new_n897));
  AOI21_X1  g696(.A(G155gat), .B1(new_n897), .B2(new_n582), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n582), .A2(G155gat), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT121), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n893), .B2(new_n900), .ZN(G1346gat));
  NAND3_X1  g700(.A1(new_n869), .A2(new_n712), .A3(new_n871), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT122), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(G162gat), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n897), .A2(new_n626), .A3(new_n692), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  OAI211_X1 g706(.A(new_n479), .B(new_n486), .C1(new_n837), .C2(new_n838), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n423), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n556), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n665), .ZN(new_n912));
  XOR2_X1   g711(.A(KEYINPUT123), .B(G176gat), .Z(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(G1349gat));
  NAND2_X1  g713(.A1(new_n909), .A2(new_n582), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n324), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n305), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n916), .B(new_n919), .C1(new_n305), .C2(new_n915), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1350gat));
  NAND2_X1  g720(.A1(new_n909), .A2(new_n692), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(G190gat), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n288), .A3(new_n712), .ZN(new_n927));
  INV_X1    g726(.A(new_n925), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n922), .A2(G190gat), .A3(new_n928), .A4(new_n923), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n684), .A2(new_n423), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n888), .A2(new_n479), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n557), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n483), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n839), .A2(new_n479), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(G197gat), .A3(new_n557), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n931), .A2(new_n479), .ZN(new_n941));
  AOI211_X1 g740(.A(new_n941), .B(new_n886), .C1(new_n887), .C2(KEYINPUT57), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n493), .B1(new_n942), .B2(new_n556), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT126), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n940), .A2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n937), .A2(G204gat), .A3(new_n666), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n889), .B2(new_n941), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n937), .A2(G204gat), .A3(new_n666), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(KEYINPUT127), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n953), .ZN(G1353gat));
  OR3_X1    g753(.A1(new_n937), .A2(G211gat), .A3(new_n763), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n942), .A2(new_n582), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n932), .B2(new_n641), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n937), .A2(G218gat), .A3(new_n729), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


