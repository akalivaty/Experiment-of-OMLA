//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT5), .ZN(new_n198));
  XNOR2_X1  g012(.A(G116), .B(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n194), .A2(new_n198), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT81), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(G104), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT85), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT82), .B1(new_n205), .B2(G104), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n211), .A3(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n206), .A3(new_n208), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT83), .B(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n205), .A2(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n204), .A2(new_n215), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n195), .A2(G116), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n200), .B(new_n202), .C1(new_n192), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n203), .A2(new_n199), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n216), .A2(new_n218), .B1(new_n223), .B2(KEYINPUT3), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n221), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT84), .B(KEYINPUT4), .Z(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n221), .A3(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G110), .B(G122), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n189), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n239), .B2(KEYINPUT87), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n244), .B(new_n226), .C1(new_n235), .C2(new_n238), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G224), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G953), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT75), .B(G125), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n256), .A3(G143), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n256), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n251), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n260), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT65), .B(G146), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G143), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n265), .B2(G143), .ZN(new_n268));
  OAI211_X1 g082(.A(KEYINPUT69), .B(new_n266), .C1(new_n268), .C2(new_n252), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(G146), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n257), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n250), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n257), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n281), .A2(KEYINPUT0), .A3(G128), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT0), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT64), .B1(new_n283), .B2(new_n252), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n262), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n252), .A3(KEYINPUT64), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n281), .B1(KEYINPUT0), .B2(G128), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n266), .A2(KEYINPUT66), .A3(new_n289), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n249), .B(new_n279), .C1(new_n286), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n248), .B1(new_n275), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n279), .B1(new_n286), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n250), .ZN(new_n294));
  INV_X1    g108(.A(new_n248), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n273), .B1(new_n263), .B2(new_n269), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n250), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n204), .A2(new_n215), .A3(new_n225), .ZN(new_n299));
  INV_X1    g113(.A(new_n238), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n233), .A2(new_n234), .ZN(new_n301));
  INV_X1    g115(.A(new_n230), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n244), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n239), .A2(KEYINPUT87), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n189), .A3(new_n306), .A4(new_n242), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n246), .A2(new_n298), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(KEYINPUT7), .B(new_n295), .C1(new_n275), .C2(new_n291), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n240), .B(KEYINPUT8), .Z(new_n310));
  NAND2_X1  g124(.A1(new_n215), .A2(new_n225), .ZN(new_n311));
  INV_X1    g125(.A(new_n204), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n313), .B2(new_n299), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n239), .B2(new_n240), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n295), .A2(KEYINPUT7), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n294), .B(new_n316), .C1(new_n296), .C2(new_n250), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n309), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G902), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n188), .B1(new_n308), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n246), .A2(new_n298), .A3(new_n307), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n187), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(KEYINPUT88), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n308), .A2(new_n320), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n187), .ZN(new_n328));
  NOR2_X1   g142(.A1(KEYINPUT96), .A2(G952), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT96), .A2(G952), .ZN(new_n331));
  AOI21_X1  g145(.A(G953), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(G234), .A2(G237), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT21), .B(G898), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(G902), .A3(G953), .A4(new_n333), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G214), .B1(G237), .B2(G902), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n325), .A2(new_n328), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n252), .A2(G143), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT13), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n259), .A2(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n342), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n206), .A2(new_n208), .ZN(new_n349));
  INV_X1    g163(.A(G122), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G116), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n191), .A2(G122), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT81), .B(G107), .ZN(new_n355));
  XNOR2_X1  g169(.A(G116), .B(G122), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n348), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n349), .A2(new_n353), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT93), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n347), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n341), .ZN(new_n363));
  XNOR2_X1  g177(.A(G128), .B(G143), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G134), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT14), .ZN(new_n367));
  OAI21_X1  g181(.A(G107), .B1(new_n352), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(new_n367), .B2(new_n356), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT9), .B(G234), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT78), .ZN(new_n372));
  INV_X1    g186(.A(G953), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G217), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n362), .A2(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n344), .B(new_n364), .ZN(new_n376));
  INV_X1    g190(.A(new_n361), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT93), .B1(new_n359), .B2(new_n360), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n372), .A2(new_n374), .ZN(new_n380));
  INV_X1    g194(.A(new_n370), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(KEYINPUT94), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n358), .A2(new_n361), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n370), .B1(new_n384), .B2(new_n376), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT94), .B1(new_n385), .B2(new_n380), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n319), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n388));
  NOR2_X1   g202(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n389));
  OAI21_X1  g203(.A(G478), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n387), .B(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n373), .A3(G214), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n259), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT68), .B(G131), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n394), .B(G143), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n250), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(G125), .A2(G140), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n249), .B2(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n253), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n405), .C1(new_n409), .C2(new_n403), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(KEYINPUT17), .A3(new_n397), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n402), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT18), .A2(G131), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n399), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n395), .A2(KEYINPUT18), .A3(G131), .ZN(new_n417));
  OAI211_X1 g231(.A(G146), .B(new_n407), .C1(new_n249), .C2(new_n404), .ZN(new_n418));
  XNOR2_X1  g232(.A(G125), .B(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n265), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT89), .B1(new_n418), .B2(new_n420), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n416), .B(new_n417), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n211), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n414), .A2(new_n426), .A3(new_n423), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n319), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  OAI21_X1  g246(.A(G475), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n419), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n265), .B(new_n435), .C1(new_n408), .C2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n401), .A2(new_n412), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n423), .A3(KEYINPUT90), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n427), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT90), .B1(new_n437), .B2(new_n423), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT91), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n423), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n427), .A4(new_n438), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n430), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n433), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n340), .A2(new_n392), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G221), .B1(new_n372), .B2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(new_n319), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n215), .A2(new_n225), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT1), .B1(new_n259), .B2(G146), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n257), .A2(new_n271), .B1(G128), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n273), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n270), .A2(new_n274), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n341), .B2(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT11), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT67), .B(new_n466), .C1(new_n341), .C2(G137), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n341), .A2(G137), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G131), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n396), .A3(new_n467), .A4(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT12), .B1(new_n463), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n273), .A2(new_n460), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n311), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n296), .B2(new_n311), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  INV_X1    g291(.A(new_n472), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n373), .A2(G227), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT80), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G140), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n458), .A2(KEYINPUT10), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n296), .A2(new_n485), .B1(new_n475), .B2(KEYINPUT10), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n293), .A2(new_n238), .A3(new_n301), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n488), .B2(new_n478), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n463), .A2(KEYINPUT12), .A3(new_n472), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n480), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n462), .A2(KEYINPUT10), .A3(new_n458), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n293), .A2(new_n238), .A3(new_n301), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT10), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n461), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n478), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n484), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n457), .B1(new_n503), .B2(new_n456), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n473), .B2(new_n479), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n484), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n489), .A2(new_n495), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(G469), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n455), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n453), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n468), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n341), .A2(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n471), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n462), .A2(KEYINPUT70), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n296), .B2(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n286), .A2(new_n290), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n472), .A3(new_n278), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n302), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n520), .B(new_n230), .C1(new_n296), .C2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n462), .A2(new_n515), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n520), .A4(new_n230), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT28), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n393), .A2(new_n373), .A3(G210), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n524), .A2(new_n527), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n520), .B(KEYINPUT30), .C1(new_n296), .C2(new_n514), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n302), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n521), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n539), .A2(new_n543), .A3(new_n536), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT29), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n531), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n525), .A2(new_n520), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n524), .B(new_n527), .C1(new_n548), .C2(new_n230), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(KEYINPUT28), .ZN(new_n550));
  INV_X1    g364(.A(new_n536), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G472), .B1(new_n546), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n521), .A2(new_n542), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n302), .A3(new_n540), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n524), .A2(new_n527), .A3(new_n536), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n532), .B2(new_n551), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n559), .A3(new_n562), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT72), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n524), .A2(new_n527), .A3(new_n536), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n543), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT72), .A3(new_n559), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  AOI211_X1 g385(.A(KEYINPUT32), .B(new_n558), .C1(new_n564), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n530), .B1(new_n538), .B2(new_n522), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n551), .B1(new_n574), .B2(new_n547), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT31), .B1(new_n543), .B2(new_n568), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT72), .B1(new_n569), .B2(new_n559), .ZN(new_n577));
  NOR4_X1   g391(.A1(new_n543), .A2(new_n568), .A3(new_n566), .A4(KEYINPUT31), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n573), .B1(new_n579), .B2(new_n557), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n556), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n411), .A2(new_n412), .ZN(new_n583));
  INV_X1    g397(.A(G110), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n252), .A2(KEYINPUT23), .A3(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n195), .A2(G128), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n195), .A2(G128), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(KEYINPUT23), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n588), .B2(KEYINPUT74), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(KEYINPUT74), .B2(new_n588), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT24), .B(G110), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT73), .ZN(new_n592));
  INV_X1    g406(.A(new_n587), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(new_n586), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT76), .B(G110), .Z(new_n597));
  OAI22_X1  g411(.A1(new_n592), .A2(new_n594), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n412), .A3(new_n420), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT22), .B(G137), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n373), .A2(G221), .A3(G234), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n599), .A3(new_n603), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n319), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT25), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT25), .A4(new_n319), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G217), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(G234), .B2(new_n319), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n605), .A2(new_n606), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(G902), .A3(new_n613), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n581), .A2(new_n582), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n582), .B1(new_n581), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n510), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(new_n222), .Z(G3));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n579), .B2(new_n319), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n558), .B1(new_n564), .B2(new_n571), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n617), .A3(new_n509), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n324), .A2(KEYINPUT98), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n187), .B1(new_n322), .B2(new_n323), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n339), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n326), .A2(KEYINPUT98), .A3(new_n187), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT99), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n630), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n321), .A2(KEYINPUT98), .A3(new_n324), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n339), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n375), .A3(new_n382), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n375), .A2(KEYINPUT33), .A3(new_n639), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(G478), .A3(new_n319), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT100), .B(G478), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n647), .B(new_n648), .C1(new_n642), .C2(new_n319), .ZN(new_n649));
  INV_X1    g463(.A(new_n648), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT101), .B1(new_n387), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n646), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT102), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n646), .B(new_n654), .C1(new_n649), .C2(new_n651), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n452), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n638), .A2(new_n337), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n628), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  OAI211_X1 g475(.A(new_n433), .B(new_n392), .C1(new_n450), .C2(new_n451), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n337), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n633), .A2(new_n663), .A3(new_n637), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n628), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND2_X1  g481(.A1(new_n611), .A2(new_n613), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n600), .B(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n319), .C1(new_n612), .C2(G234), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n509), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n626), .A3(new_n453), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AND2_X1   g490(.A1(new_n581), .A2(new_n673), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n373), .A2(G900), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n333), .A2(G902), .ZN(new_n680));
  OR3_X1    g494(.A1(new_n679), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n334), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n638), .A2(new_n662), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT104), .B(G128), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G30));
  AND2_X1   g502(.A1(new_n452), .A2(new_n392), .ZN(new_n689));
  INV_X1    g503(.A(new_n672), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n339), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT106), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n683), .B(KEYINPUT39), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n509), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n325), .A2(new_n328), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n692), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n551), .B1(new_n561), .B2(new_n538), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n319), .B1(new_n549), .B2(new_n536), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n572), .B2(new_n580), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n698), .B(new_n705), .C1(KEYINPUT40), .C2(new_n694), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR2_X1   g521(.A1(new_n638), .A2(new_n657), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n677), .A2(new_n708), .A3(new_n683), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  INV_X1    g524(.A(new_n484), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n500), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n490), .A2(new_n491), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(KEYINPUT86), .B2(new_n713), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n714), .A2(new_n493), .B1(new_n484), .B2(new_n501), .ZN(new_n715));
  OAI211_X1 g529(.A(KEYINPUT107), .B(G469), .C1(new_n715), .C2(G902), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n503), .B2(new_n456), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n494), .A2(new_n502), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n456), .A3(new_n319), .ZN(new_n721));
  INV_X1    g535(.A(new_n455), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n719), .A2(new_n724), .A3(new_n617), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n658), .A2(new_n581), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n664), .A2(new_n581), .A3(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AND2_X1   g544(.A1(new_n633), .A2(new_n637), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n723), .B1(new_n718), .B2(new_n716), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n690), .A2(new_n452), .A3(new_n392), .A4(new_n337), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n581), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  INV_X1    g549(.A(new_n732), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n638), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n581), .A4(new_n733), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT109), .B(G119), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G21));
  OAI21_X1  g556(.A(new_n576), .B1(new_n550), .B2(new_n536), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n558), .B1(new_n744), .B2(new_n571), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n624), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n725), .A2(new_n746), .A3(new_n338), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n633), .A2(new_n637), .A3(new_n689), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n350), .ZN(G24));
  NOR2_X1   g564(.A1(new_n577), .A2(new_n578), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n557), .B1(new_n751), .B2(new_n743), .ZN(new_n752));
  AOI21_X1  g566(.A(G902), .B1(new_n564), .B2(new_n571), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n752), .B(new_n672), .C1(new_n753), .C2(new_n623), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n656), .A2(new_n452), .A3(new_n683), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n547), .B1(new_n528), .B2(KEYINPUT28), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n551), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n552), .B1(new_n761), .B2(new_n544), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n623), .B1(new_n762), .B2(new_n554), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n576), .B1(new_n760), .B2(new_n536), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n557), .B1(new_n751), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT32), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n579), .A2(new_n573), .A3(new_n557), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n617), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n759), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n581), .A2(KEYINPUT111), .A3(new_n617), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n656), .A2(new_n452), .A3(new_n683), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n505), .A2(new_n484), .B1(new_n489), .B2(new_n495), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(G469), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n711), .B1(new_n713), .B2(new_n500), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n495), .A2(new_n500), .A3(new_n711), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT110), .A4(new_n456), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n455), .B1(new_n779), .B2(new_n504), .ZN(new_n780));
  INV_X1    g594(.A(new_n339), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n325), .B2(new_n328), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT42), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n770), .A2(new_n771), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n508), .A2(KEYINPUT110), .ZN(new_n787));
  INV_X1    g601(.A(new_n457), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n774), .A2(new_n773), .A3(G469), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n721), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n782), .A2(new_n722), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n581), .A2(new_n617), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n784), .B1(new_n793), .B2(new_n755), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NOR2_X1   g610(.A1(new_n662), .A2(new_n684), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n581), .A2(new_n617), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  INV_X1    g613(.A(new_n656), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n452), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n800), .A2(KEYINPUT43), .A3(new_n452), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n626), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n672), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n774), .A2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n774), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT46), .B1(new_n813), .B2(new_n788), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n456), .B2(new_n503), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n455), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n693), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n782), .B(KEYINPUT113), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n807), .B2(new_n808), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n810), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NAND2_X1  g638(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n817), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n768), .A2(new_n769), .A3(new_n772), .A4(new_n782), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(new_n404), .ZN(G42));
  INV_X1    g645(.A(new_n748), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n672), .A2(new_n684), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n702), .A3(new_n780), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n709), .A2(new_n686), .A3(new_n757), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n677), .A2(new_n685), .B1(new_n756), .B2(new_n737), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n709), .A4(new_n834), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n729), .A2(new_n674), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n340), .B1(new_n662), .B2(new_n657), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n626), .A2(new_n842), .A3(new_n617), .A4(new_n509), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n747), .B2(new_n748), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n740), .A3(new_n621), .A4(new_n726), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n791), .A2(new_n755), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n624), .A2(new_n690), .A3(new_n745), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT115), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n783), .A2(new_n754), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n452), .A2(new_n392), .A3(new_n684), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n581), .A2(new_n673), .A3(new_n782), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n798), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n795), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT116), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n798), .B(new_n854), .C1(new_n849), .C2(new_n851), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n786), .B2(new_n794), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  INV_X1    g675(.A(new_n726), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n841), .A3(new_n844), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT77), .B1(new_n768), .B2(new_n769), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n618), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n865), .A2(new_n510), .B1(new_n735), .B2(new_n739), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n860), .A2(new_n861), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n840), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT53), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n837), .A2(new_n838), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n871), .B(new_n840), .C1(new_n858), .C2(new_n867), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n836), .A2(new_n839), .ZN(new_n875));
  INV_X1    g689(.A(new_n846), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n860), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n874), .B(new_n879), .C1(new_n868), .C2(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n732), .A2(new_n782), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n769), .A3(new_n334), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n703), .A2(new_n704), .A3(new_n883), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n884), .A2(new_n452), .A3(new_n656), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n803), .A2(new_n882), .A3(new_n334), .A4(new_n804), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n848), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n769), .A2(new_n334), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n805), .A2(new_n746), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n697), .A2(new_n339), .A3(new_n736), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT50), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n885), .B(new_n887), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n719), .A2(new_n455), .A3(new_n721), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n821), .B(new_n889), .C1(new_n828), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  OR3_X1    g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n332), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n884), .A2(new_n657), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n899), .B(new_n900), .C1(new_n737), .C2(new_n890), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n770), .A2(new_n771), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n886), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n901), .B2(KEYINPUT117), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n898), .A2(new_n902), .A3(new_n903), .A4(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n881), .A2(new_n909), .B1(G952), .B2(G953), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n719), .A2(new_n721), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(KEYINPUT49), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n769), .A2(new_n455), .A3(new_n781), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n801), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(KEYINPUT49), .ZN(new_n915));
  OR4_X1    g729(.A1(new_n697), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n705), .B2(new_n916), .ZN(G75));
  OAI21_X1  g731(.A(new_n879), .B1(new_n868), .B2(KEYINPUT53), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G210), .A3(G902), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n246), .A2(new_n307), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n298), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n308), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT119), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n919), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n919), .B2(new_n920), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n373), .A2(G952), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT120), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n880), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n457), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n720), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n813), .B(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n918), .A2(G902), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n928), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n918), .A2(G902), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n447), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n928), .ZN(G60));
  NAND2_X1  g761(.A1(new_n644), .A2(new_n645), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT59), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n933), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n929), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n949), .B1(new_n881), .B2(new_n951), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G63));
  XNOR2_X1  g770(.A(new_n615), .B(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n918), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n930), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n918), .A2(new_n670), .A3(new_n961), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n962), .A3(new_n930), .ZN(new_n967));
  XNOR2_X1  g781(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G66));
  OAI21_X1  g783(.A(G953), .B1(new_n335), .B2(new_n247), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n876), .B2(G953), .ZN(new_n971));
  INV_X1    g785(.A(G898), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n921), .B1(new_n972), .B2(G953), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n971), .B(new_n973), .Z(G69));
  NAND2_X1  g788(.A1(new_n560), .A2(new_n540), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n435), .B1(new_n408), .B2(new_n434), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT126), .Z(new_n977));
  XOR2_X1   g791(.A(new_n975), .B(new_n977), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n837), .A2(new_n709), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n706), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n706), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  INV_X1    g798(.A(new_n782), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n985), .B(new_n694), .C1(new_n657), .C2(new_n662), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n830), .B1(new_n865), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n823), .A2(new_n982), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n979), .B1(new_n988), .B2(new_n373), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n823), .A2(new_n795), .ZN(new_n990));
  INV_X1    g804(.A(new_n830), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n819), .A2(new_n904), .A3(new_n832), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n798), .A3(new_n980), .A4(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n373), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n679), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n989), .B1(new_n995), .B2(new_n979), .ZN(new_n996));
  NAND2_X1  g810(.A1(G227), .A2(G900), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(G953), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G72));
  NOR3_X1   g813(.A1(new_n990), .A2(new_n846), .A3(new_n993), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n544), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n988), .B2(new_n846), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n699), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1004), .B(new_n1006), .C1(G952), .C2(new_n373), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n869), .A2(new_n872), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n544), .A2(new_n699), .A3(new_n1003), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(G57));
endmodule


