//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G77), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT9), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n215), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n253), .A2(new_n255), .B1(G150), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n215), .A3(new_n247), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n261), .A2(new_n263), .B1(G50), .B2(new_n260), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(new_n266), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n246), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n269), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(G223), .B1(new_n279), .B2(new_n218), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G222), .A3(new_n273), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n289), .A3(G274), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n286), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(G226), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT66), .B(G200), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G190), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n270), .A2(new_n272), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n270), .A2(new_n272), .A3(new_n302), .A4(new_n300), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n304), .B2(new_n303), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n253), .A2(new_n262), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n308), .A2(new_n261), .B1(new_n260), .B2(new_n253), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n274), .A2(new_n207), .A3(new_n275), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT7), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT7), .B1(new_n279), .B2(new_n207), .ZN(new_n315));
  OAI21_X1  g0115(.A(G68), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G68), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n202), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G58), .A2(G68), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n256), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n249), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(KEYINPUT16), .A3(new_n323), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n311), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G274), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n284), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(G232), .A2(new_n293), .B1(new_n330), .B2(new_n287), .ZN(new_n331));
  OAI211_X1 g0131(.A(G223), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n332));
  OAI211_X1 g0132(.A(G226), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n333));
  INV_X1    g0133(.A(G87), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n254), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n284), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n331), .A2(new_n336), .A3(G179), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT18), .B1(new_n328), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n331), .A2(new_n336), .A3(G190), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n312), .A2(new_n313), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n317), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n325), .B1(new_n347), .B2(new_n322), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n327), .A2(new_n348), .A3(new_n248), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n309), .B(KEYINPUT75), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n338), .A2(new_n339), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n349), .A2(new_n350), .A3(new_n343), .A4(new_n342), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n341), .A2(new_n351), .A3(new_n355), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n295), .A2(G179), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n265), .B(new_n361), .C1(new_n362), .C2(new_n295), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n276), .A2(G238), .B1(new_n279), .B2(G107), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n281), .A2(G232), .A3(new_n273), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n284), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n291), .B1(G244), .B2(new_n293), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n297), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n255), .B1(new_n218), .B2(G20), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n253), .A2(new_n256), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n249), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n262), .A2(G77), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n261), .A2(new_n377), .B1(new_n218), .B2(new_n260), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n371), .B(new_n379), .C1(new_n380), .C2(new_n370), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n370), .B2(new_n362), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n368), .A2(new_n383), .A3(new_n369), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n307), .A2(new_n360), .A3(new_n364), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n260), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n317), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT12), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n255), .A2(G77), .B1(G20), .B2(new_n317), .ZN(new_n391));
  INV_X1    g0191(.A(new_n256), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n201), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n394));
  INV_X1    g0194(.A(new_n261), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(G68), .A3(new_n262), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT11), .B1(new_n393), .B2(new_n248), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT69), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n281), .A2(KEYINPUT69), .A3(G226), .A4(new_n273), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n281), .A2(G232), .A3(G1698), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n284), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n290), .B1(new_n410), .B2(new_n292), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n401), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(KEYINPUT13), .B(new_n411), .C1(new_n408), .C2(new_n284), .ZN(new_n414));
  OAI21_X1  g0214(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT14), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(new_n401), .A3(new_n412), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n409), .A2(new_n412), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n401), .A4(new_n412), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n422), .A2(new_n424), .A3(G179), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(G169), .C1(new_n413), .C2(new_n414), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n400), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n362), .B1(new_n424), .B2(new_n420), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT73), .B1(new_n431), .B2(new_n427), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT14), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n429), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(KEYINPUT74), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n399), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n422), .A2(new_n424), .A3(G190), .A4(new_n425), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n438), .A2(new_n399), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n413), .B2(new_n414), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT70), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT70), .B(G200), .C1(new_n413), .C2(new_n414), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n439), .A2(new_n444), .A3(KEYINPUT72), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT72), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n387), .A2(new_n437), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n206), .A2(G33), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n249), .A2(new_n260), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT25), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n260), .B2(G107), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n260), .A2(new_n452), .A3(G107), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n451), .A2(G107), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n207), .B(G87), .C1(new_n277), .C2(new_n278), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n281), .A2(new_n460), .A3(new_n207), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT23), .ZN(new_n465));
  INV_X1    g0265(.A(G107), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n468), .A2(KEYINPUT81), .B1(new_n469), .B2(G20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT24), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n457), .B1(new_n473), .B2(new_n248), .ZN(new_n474));
  OAI211_X1 g0274(.A(G250), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT82), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n276), .B2(G257), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n284), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(KEYINPUT83), .A3(new_n284), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  INV_X1    g0289(.A(new_n215), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n487), .A2(new_n489), .B1(new_n490), .B2(new_n288), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n206), .A2(G45), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G274), .A3(new_n289), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n485), .A2(new_n486), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G169), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n493), .B1(new_n482), .B2(new_n284), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G179), .A3(new_n499), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n474), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n472), .A2(KEYINPUT24), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n462), .B2(new_n471), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n248), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n456), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n485), .A2(new_n380), .A3(new_n486), .A4(new_n501), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n475), .A2(new_n476), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n276), .A2(new_n478), .A3(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n499), .B(new_n492), .C1(new_n516), .C2(new_n289), .ZN(new_n517));
  INV_X1    g0317(.A(G200), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n506), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n273), .B(new_n522), .C1(new_n277), .C2(new_n278), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n220), .B1(new_n274), .B2(new_n275), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g0326(.A(G250), .B1(new_n277), .B2(new_n278), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n273), .B1(new_n527), .B2(KEYINPUT4), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n284), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n497), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n489), .B1(new_n530), .B2(new_n495), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G257), .A3(new_n289), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n499), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n533), .A3(new_n383), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n499), .A2(new_n532), .ZN(new_n535));
  INV_X1    g0335(.A(G250), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n274), .B2(new_n275), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(G1698), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G244), .B1(new_n277), .B2(new_n278), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n538), .B1(G33), .B2(G283), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n541), .A3(new_n523), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n535), .B1(new_n542), .B2(new_n284), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n534), .B1(new_n543), .B2(G169), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n260), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n450), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT76), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  AND2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n466), .A2(KEYINPUT6), .A3(G97), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n207), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G77), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n392), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n549), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(G107), .B1(new_n314), .B2(new_n315), .ZN(new_n559));
  INV_X1    g0359(.A(new_n557), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n466), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n550), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT76), .B(new_n560), .C1(new_n563), .C2(new_n207), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n548), .B1(new_n565), .B2(new_n248), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n544), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n248), .ZN(new_n568));
  INV_X1    g0368(.A(new_n548), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n529), .A2(new_n533), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n380), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT77), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n518), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n574), .B2(new_n571), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n567), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n491), .A2(G270), .B1(new_n330), .B2(new_n498), .ZN(new_n578));
  OAI211_X1 g0378(.A(G257), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n579));
  OAI211_X1 g0379(.A(G264), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n274), .A2(G303), .A3(new_n275), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n284), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n583), .A3(G179), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n247), .A2(new_n215), .B1(G20), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n524), .B(new_n207), .C1(G33), .C2(new_n547), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n388), .A2(new_n587), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n587), .C2(new_n450), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n450), .B2(new_n587), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n593), .B2(new_n592), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT79), .B1(new_n599), .B2(new_n584), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n578), .A2(new_n583), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n596), .A2(G169), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(KEYINPUT80), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(KEYINPUT80), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n596), .A2(new_n602), .A3(G169), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(G200), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(new_n599), .C1(new_n380), .C2(new_n602), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n601), .A2(new_n605), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n450), .A2(new_n372), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n373), .A2(new_n260), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n281), .A2(new_n207), .A3(G68), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n552), .A2(new_n334), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n406), .A2(new_n207), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n254), .A2(new_n547), .A3(KEYINPUT19), .A4(G20), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT78), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n249), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n613), .B(KEYINPUT78), .C1(new_n617), .C2(new_n618), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n611), .B(new_n612), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n536), .B1(new_n488), .B2(G1), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n206), .A2(new_n329), .A3(G45), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n289), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(G238), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G33), .A2(G116), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n540), .C2(new_n273), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n284), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n383), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G169), .B2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(G190), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n296), .B2(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(new_n612), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n450), .A2(new_n334), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n639));
  AOI21_X1  g0439(.A(G20), .B1(G33), .B2(G97), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT19), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n255), .A2(new_n614), .A3(G97), .ZN(new_n642));
  AOI21_X1  g0442(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(G68), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n248), .B1(new_n644), .B2(KEYINPUT78), .ZN(new_n645));
  INV_X1    g0445(.A(new_n622), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n636), .B(new_n638), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n623), .A2(new_n633), .B1(new_n635), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n610), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n448), .A2(new_n521), .A3(new_n577), .A4(new_n649), .ZN(G372));
  XNOR2_X1  g0450(.A(new_n626), .B(KEYINPUT84), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n630), .A2(new_n284), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n362), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(KEYINPUT85), .A3(new_n632), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT85), .ZN(new_n656));
  AOI21_X1  g0456(.A(G169), .B1(new_n651), .B2(new_n652), .ZN(new_n657));
  AOI211_X1 g0457(.A(G179), .B(new_n627), .C1(new_n630), .C2(new_n284), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n623), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n635), .A2(new_n647), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n567), .C1(new_n623), .C2(new_n633), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n529), .A2(new_n533), .A3(new_n383), .ZN(new_n664));
  AOI21_X1  g0464(.A(G169), .B1(new_n529), .B2(new_n533), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT86), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n570), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT86), .B1(new_n544), .B2(new_n566), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n653), .A2(new_n297), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n634), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n647), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n512), .A2(new_n519), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n474), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n577), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n601), .A2(new_n605), .A3(new_n607), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n506), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n663), .B(new_n676), .C1(new_n679), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n448), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n351), .A2(new_n358), .ZN(new_n684));
  INV_X1    g0484(.A(new_n399), .ZN(new_n685));
  AOI211_X1 g0485(.A(new_n400), .B(new_n429), .C1(new_n432), .C2(new_n433), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT74), .B1(new_n434), .B2(new_n435), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n385), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n445), .B2(new_n446), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n684), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n341), .A2(new_n355), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n307), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n683), .A2(new_n364), .A3(new_n693), .ZN(G369));
  NAND3_X1  g0494(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n511), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT87), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n521), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT88), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n702), .A4(new_n703), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n506), .A2(new_n700), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n700), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n599), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n680), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n610), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n680), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n700), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n706), .A2(new_n707), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n506), .A2(new_n711), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n716), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n210), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n615), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n213), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n671), .B1(new_n670), .B2(new_n675), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n636), .B1(new_n372), .B2(new_n450), .C1(new_n645), .C2(new_n646), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT85), .B1(new_n654), .B2(new_n632), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n657), .A2(new_n658), .A3(new_n656), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT91), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n577), .A2(new_n675), .A3(new_n678), .ZN(new_n738));
  INV_X1    g0538(.A(new_n506), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n717), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n647), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n634), .A3(new_n672), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n735), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n668), .A2(new_n669), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT26), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n666), .A2(new_n570), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n648), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n660), .B1(new_n748), .B2(new_n671), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT91), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n737), .A2(new_n741), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n730), .B1(new_n752), .B2(new_n711), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n682), .A2(new_n711), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(KEYINPUT29), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(G179), .B1(new_n578), .B2(new_n583), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(new_n653), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT89), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(new_n517), .A4(new_n571), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n504), .A2(new_n543), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n631), .A2(G179), .A3(new_n583), .A4(new_n578), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n517), .A2(new_n571), .A3(new_n757), .A4(new_n653), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT89), .ZN(new_n766));
  INV_X1    g0566(.A(new_n763), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n767), .A2(KEYINPUT30), .A3(new_n504), .A4(new_n543), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n760), .A2(new_n764), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n700), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT90), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n521), .A2(new_n649), .A3(new_n577), .A4(new_n711), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n764), .A2(new_n768), .A3(new_n765), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT90), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n770), .A2(new_n777), .A3(new_n771), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n773), .A2(new_n774), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G330), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n729), .B1(new_n782), .B2(G1), .ZN(G364));
  NAND2_X1  g0583(.A1(new_n207), .A2(G13), .ZN(new_n784));
  OAI21_X1  g0584(.A(G1), .B1(new_n784), .B2(new_n488), .ZN(new_n785));
  OR3_X1    g0585(.A1(new_n724), .A2(KEYINPUT93), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT93), .B1(new_n724), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n723), .A2(new_n281), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n488), .B2(new_n214), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n241), .B2(new_n488), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n210), .A2(new_n281), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT94), .Z(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n587), .B2(new_n723), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OR3_X1    g0596(.A1(KEYINPUT95), .A2(G13), .A3(G33), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT95), .B1(G13), .B2(G33), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n215), .B1(G20), .B2(new_n362), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n788), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT96), .ZN(new_n805));
  INV_X1    g0605(.A(new_n801), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n297), .A2(G20), .A3(new_n383), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G190), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n380), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n807), .A2(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n207), .A2(new_n383), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(G200), .B1(new_n816), .B2(KEYINPUT97), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(KEYINPUT97), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G190), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G311), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n380), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G322), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G179), .A2(G200), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G190), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n281), .B1(new_n825), .B2(G294), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n816), .A2(new_n380), .A3(new_n518), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n816), .A2(G190), .A3(new_n518), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G326), .A2(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n820), .A2(new_n822), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n823), .A2(G20), .A3(new_n380), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT98), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT98), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n814), .B(new_n831), .C1(G329), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(KEYINPUT99), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(KEYINPUT99), .ZN(new_n841));
  INV_X1    g0641(.A(G159), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT32), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n281), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n812), .A2(new_n334), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G107), .C2(new_n809), .ZN(new_n847));
  INV_X1    g0647(.A(new_n825), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n547), .ZN(new_n849));
  INV_X1    g0649(.A(new_n828), .ZN(new_n850));
  INV_X1    g0650(.A(new_n827), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n850), .A2(new_n317), .B1(new_n851), .B2(new_n201), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n849), .B(new_n852), .C1(new_n844), .C2(new_n843), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n819), .A2(new_n218), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n821), .A2(G58), .ZN(new_n855));
  AND4_X1   g0655(.A1(new_n847), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n840), .A2(new_n841), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n802), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n805), .B1(new_n714), .B2(new_n806), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT100), .Z(new_n860));
  XOR2_X1   g0660(.A(new_n715), .B(KEYINPUT92), .Z(new_n861));
  OAI21_X1  g0661(.A(new_n788), .B1(new_n714), .B2(G330), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(G396));
  INV_X1    g0663(.A(new_n788), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n381), .B1(new_n379), .B2(new_n711), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n385), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n689), .A2(new_n711), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n754), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n682), .A2(new_n868), .A3(new_n711), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n864), .B1(new_n872), .B2(new_n780), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n780), .B2(new_n872), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G137), .A2(new_n827), .B1(new_n828), .B2(G150), .ZN(new_n875));
  INV_X1    g0675(.A(new_n819), .ZN(new_n876));
  INV_X1    g0676(.A(new_n821), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT101), .B(G143), .Z(new_n878));
  OAI221_X1 g0678(.A(new_n875), .B1(new_n876), .B2(new_n842), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT34), .Z(new_n880));
  AOI22_X1  g0680(.A1(new_n837), .A2(G132), .B1(G50), .B2(new_n811), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n809), .A2(G68), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n279), .B1(new_n825), .B2(G58), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n809), .A2(G87), .ZN(new_n885));
  INV_X1    g0685(.A(G311), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n885), .B1(new_n836), .B2(new_n886), .C1(new_n812), .C2(new_n466), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n850), .A2(new_n807), .B1(new_n851), .B2(new_n813), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n281), .B(new_n888), .C1(G97), .C2(new_n825), .ZN(new_n889));
  INV_X1    g0689(.A(G294), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n889), .B1(new_n876), .B2(new_n587), .C1(new_n890), .C2(new_n877), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n880), .A2(new_n884), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n802), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n799), .A2(new_n802), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n788), .B1(new_n556), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n895), .C1(new_n868), .C2(new_n800), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n874), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(G384));
  INV_X1    g0698(.A(new_n563), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(G116), .A4(new_n216), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT36), .Z(new_n903));
  OAI211_X1 g0703(.A(new_n218), .B(new_n214), .C1(new_n202), .C2(new_n317), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n201), .A2(G68), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n206), .B(G13), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n871), .A2(new_n867), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n399), .A2(new_n711), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n437), .A2(new_n447), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n909), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n445), .A2(new_n446), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n688), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n309), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n698), .B1(new_n349), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n359), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n352), .A2(new_n354), .ZN(new_n918));
  INV_X1    g0718(.A(new_n698), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n352), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(new_n356), .ZN(new_n922));
  AND4_X1   g0722(.A1(new_n349), .A2(new_n350), .A3(new_n343), .A4(new_n342), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n349), .A2(new_n915), .B1(new_n338), .B2(new_n339), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(new_n916), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(new_n925), .B2(new_n921), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n917), .A2(new_n926), .A3(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n917), .A2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n914), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n692), .A2(new_n698), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n917), .A2(new_n926), .A3(KEYINPUT38), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n918), .A2(new_n920), .A3(new_n356), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT37), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n922), .ZN(new_n937));
  INV_X1    g0737(.A(new_n920), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n359), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n933), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n437), .A2(new_n711), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n932), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n931), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n448), .B1(new_n753), .B2(new_n755), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n947), .A2(new_n364), .A3(new_n693), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n946), .B(new_n948), .Z(new_n949));
  NAND3_X1  g0749(.A1(new_n769), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n774), .A2(new_n950), .A3(new_n772), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n448), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT102), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n430), .A2(new_n436), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n685), .B(new_n700), .C1(new_n954), .C2(new_n447), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n688), .A2(new_n912), .A3(new_n911), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n934), .A2(new_n940), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n951), .A2(new_n868), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT40), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT40), .B1(new_n930), .B2(new_n927), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n957), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n953), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n953), .A2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(G330), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n949), .A2(new_n968), .B1(G1), .B2(new_n784), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT103), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n969), .A2(new_n970), .B1(new_n949), .B2(new_n968), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n907), .B1(new_n971), .B2(new_n972), .ZN(G367));
  AOI211_X1 g0773(.A(new_n802), .B(new_n801), .C1(new_n723), .C2(new_n373), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n789), .A2(new_n236), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n788), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n742), .A2(new_n711), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n660), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n744), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n279), .B1(new_n832), .B2(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n851), .A2(new_n886), .B1(new_n466), .B2(new_n848), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(G294), .C2(new_n828), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n811), .A2(G116), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT46), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n809), .A2(G97), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G283), .A2(new_n819), .B1(new_n821), .B2(G303), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n279), .B1(new_n809), .B2(new_n218), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n825), .A2(G68), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n851), .B2(new_n878), .C1(new_n842), .C2(new_n850), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G150), .B2(new_n821), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n990), .B(new_n993), .C1(new_n201), .C2(new_n876), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n811), .A2(G58), .B1(G137), .B2(new_n833), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT108), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n988), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT109), .Z(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n976), .B1(new_n806), .B2(new_n979), .C1(new_n999), .C2(new_n858), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n724), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n719), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n718), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(new_n710), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n861), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n708), .A2(new_n709), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n719), .B1(new_n1006), .B2(new_n718), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n715), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1005), .A2(new_n781), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n570), .A2(new_n700), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n577), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n567), .A2(new_n700), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT104), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT104), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1015), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n719), .A2(new_n1017), .A3(new_n720), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT45), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT44), .B1(new_n721), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1022), .B(new_n1017), .C1(new_n719), .C2(new_n720), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n716), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1018), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n716), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1009), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1001), .B1(new_n1030), .B2(new_n782), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n785), .B(KEYINPUT106), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n719), .A2(new_n1020), .A3(KEYINPUT42), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n747), .B1(new_n1020), .B2(new_n739), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n711), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT42), .B1(new_n719), .B2(new_n1020), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n979), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1002), .A2(new_n1017), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(KEYINPUT42), .B1(new_n1035), .B2(new_n711), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1045), .A2(new_n1040), .A3(new_n1039), .A4(new_n1034), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1028), .B2(new_n1020), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1028), .A2(new_n1020), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1043), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT105), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT105), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1043), .A2(new_n1046), .A3(new_n1052), .A4(new_n1049), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1000), .B1(new_n1033), .B2(new_n1054), .ZN(G387));
  NOR2_X1   g0855(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n1032), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n812), .A2(new_n219), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G150), .B2(new_n833), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT110), .Z(new_n1060));
  NOR2_X1   g0860(.A1(new_n848), .A2(new_n372), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n253), .B2(new_n828), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n279), .B1(new_n827), .B2(G159), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1062), .A2(new_n986), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G50), .A2(new_n821), .B1(new_n819), .B2(G68), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n281), .B1(new_n833), .B2(G326), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n812), .A2(new_n890), .B1(new_n807), .B2(new_n848), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G322), .A2(new_n827), .B1(new_n828), .B2(G311), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n876), .B2(new_n813), .C1(new_n980), .C2(new_n877), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT49), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1067), .B1(new_n587), .B2(new_n810), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1066), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n802), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n233), .A2(new_n488), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n726), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1079), .A2(new_n789), .B1(new_n1080), .B2(new_n794), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n253), .A2(new_n201), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT50), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n488), .B1(new_n317), .B2(new_n556), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1083), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1081), .A2(new_n1085), .B1(G107), .B2(new_n210), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n788), .B1(new_n1086), .B2(new_n803), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1078), .B(new_n1087), .C1(new_n1006), .C2(new_n806), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1009), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n724), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1056), .A2(new_n782), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1057), .B(new_n1088), .C1(new_n1090), .C2(new_n1091), .ZN(G393));
  NAND3_X1  g0892(.A1(new_n1025), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n803), .B1(new_n547), .B2(new_n210), .C1(new_n790), .C2(new_n244), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n864), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n828), .A2(G50), .B1(new_n825), .B2(G77), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n253), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n876), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT111), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n821), .A2(G159), .B1(G150), .B2(new_n827), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  OAI211_X1 g0901(.A(new_n885), .B(new_n281), .C1(new_n832), .C2(new_n878), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G68), .B2(new_n811), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n821), .A2(G311), .B1(G317), .B2(new_n827), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT113), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n281), .B1(new_n833), .B2(G322), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n850), .B2(new_n813), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n825), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G107), .A2(new_n809), .B1(new_n811), .B2(G283), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n890), .C2(new_n876), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1104), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1095), .B1(new_n1114), .B2(new_n802), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1017), .B2(new_n806), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1093), .A2(KEYINPUT114), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1089), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n724), .A3(new_n1030), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(G390));
  NAND3_X1  g0925(.A1(new_n951), .A2(G330), .A3(new_n868), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n956), .B2(new_n955), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n941), .A2(new_n942), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n914), .B2(new_n944), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n958), .A2(new_n944), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n752), .A2(new_n711), .A3(new_n866), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n867), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1132), .B2(new_n957), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1127), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n779), .A2(G330), .A3(new_n868), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1135), .A2(new_n956), .A3(new_n955), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n908), .B1(new_n1136), .B2(new_n1127), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n780), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n957), .A2(new_n1138), .A3(new_n868), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n867), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n746), .A2(new_n749), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(KEYINPUT91), .B1(new_n738), .B2(new_n740), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n700), .B1(new_n1142), .B2(new_n751), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1143), .B2(new_n866), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1126), .A2(new_n955), .A3(new_n956), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1130), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n910), .A2(new_n913), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n955), .A2(new_n956), .B1(new_n867), .B2(new_n871), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n944), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n943), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1153), .A3(new_n1139), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n448), .A2(G330), .A3(new_n951), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n364), .A2(new_n947), .A3(new_n1155), .A4(new_n693), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1134), .A2(new_n1147), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n724), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT115), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1158), .A2(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(KEYINPUT115), .A3(new_n724), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1128), .A2(new_n800), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n894), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n828), .A2(G137), .B1(new_n825), .B2(G159), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n876), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT117), .Z(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n281), .B1(new_n1171), .B2(new_n851), .C1(new_n836), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G50), .B2(new_n809), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n811), .A2(G150), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT53), .Z(new_n1176));
  INV_X1    g0976(.A(G132), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1174), .B(new_n1176), .C1(new_n1177), .C2(new_n877), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT118), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT118), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n281), .B1(new_n825), .B2(G77), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G283), .A2(new_n827), .B1(new_n828), .B2(G107), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n877), .C2(new_n587), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G97), .B2(new_n819), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n846), .B1(G68), .B2(new_n809), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n890), .C2(new_n836), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1180), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n864), .B1(new_n253), .B2(new_n1166), .C1(new_n1188), .C2(new_n858), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1165), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT116), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1032), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1161), .B2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1134), .A2(new_n1154), .A3(KEYINPUT116), .A4(new_n1032), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1164), .A2(new_n1195), .ZN(G378));
  AND2_X1   g0996(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1156), .B1(new_n1161), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT121), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1157), .A2(KEYINPUT121), .A3(new_n1156), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n307), .A2(new_n364), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n698), .B1(new_n271), .B2(new_n267), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR3_X1    g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n957), .A2(new_n959), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1213), .A2(new_n962), .B1(new_n960), .B2(KEYINPUT40), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1214), .B2(new_n967), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n964), .A2(G330), .A3(new_n1211), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n946), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n946), .A3(new_n1216), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1202), .A2(KEYINPUT57), .A3(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1157), .A2(KEYINPUT121), .A3(new_n1156), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT121), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1219), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n1217), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n724), .B(new_n1221), .C1(new_n1227), .C2(KEYINPUT57), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n812), .A2(new_n1168), .B1(new_n1177), .B2(new_n850), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G137), .B2(new_n819), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1171), .B2(new_n877), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n827), .A2(G125), .B1(new_n825), .B2(G150), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT119), .Z(new_n1233));
  NOR2_X1   g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1237));
  INV_X1    g1037(.A(G41), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(KEYINPUT120), .B(G124), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n254), .B(new_n1238), .C1(new_n1239), .C2(new_n832), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n809), .B2(G159), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1236), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G116), .A2(new_n827), .B1(new_n828), .B2(G97), .ZN(new_n1243));
  AND4_X1   g1043(.A1(new_n1238), .A2(new_n1243), .A3(new_n279), .A4(new_n991), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n466), .B2(new_n877), .C1(new_n372), .C2(new_n876), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n836), .A2(new_n807), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n810), .A2(new_n202), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1245), .A2(new_n1058), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT58), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G50), .B1(new_n254), .B2(new_n1238), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n281), .B2(G41), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1248), .A2(KEYINPUT58), .ZN(new_n1252));
  AND4_X1   g1052(.A1(new_n1242), .A2(new_n1249), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n864), .B1(G50), .B2(new_n1166), .C1(new_n1253), .C2(new_n858), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1212), .B2(new_n799), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1220), .B2(new_n1032), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1228), .A2(new_n1256), .ZN(G375));
  INV_X1    g1057(.A(new_n1156), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1197), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1001), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1160), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT122), .Z(new_n1262));
  AOI21_X1  g1062(.A(new_n788), .B1(new_n317), .B2(new_n894), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT124), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G294), .A2(new_n827), .B1(new_n828), .B2(G116), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n876), .B2(new_n466), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT125), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n281), .B(new_n1061), .C1(new_n837), .C2(G303), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G77), .A2(new_n809), .B1(new_n811), .B2(G97), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n807), .C2(new_n877), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n281), .B1(new_n851), .B2(new_n1177), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n850), .A2(new_n1168), .B1(new_n201), .B2(new_n848), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1271), .B(new_n1272), .C1(G137), .C2(new_n821), .ZN(new_n1273));
  INV_X1    g1073(.A(G150), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n876), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1247), .B1(G128), .B2(new_n837), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n842), .B2(new_n812), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1267), .A2(new_n1270), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1264), .B1(new_n1278), .B2(new_n802), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n957), .B2(new_n800), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1032), .B(KEYINPUT123), .Z(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1197), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1262), .A2(new_n1283), .ZN(G381));
  AND3_X1   g1084(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1000), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1287));
  OR2_X1    g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(G381), .A2(new_n1287), .A3(G384), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1195), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1289), .A2(new_n1291), .A3(new_n1228), .A4(new_n1256), .ZN(G407));
  NAND2_X1  g1092(.A1(new_n699), .A2(G213), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G407), .B(G213), .C1(G375), .C2(new_n1295), .ZN(G409));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(G387), .A2(G390), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1286), .A2(new_n1000), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G387), .A2(G390), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1287), .A3(new_n1297), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1217), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n724), .B1(new_n1224), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1220), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G378), .B(new_n1256), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1260), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1226), .B1(new_n1309), .B2(new_n1281), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1291), .B1(new_n1310), .B2(new_n1255), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1293), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1294), .A2(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1259), .B(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1160), .A2(new_n724), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1319), .B2(new_n1283), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n897), .B(new_n1282), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1315), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1259), .B(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(new_n1317), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n897), .B1(new_n1325), .B2(new_n1282), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1319), .A2(G384), .A3(new_n1283), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1314), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1322), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1312), .A2(new_n1293), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1304), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1312), .A2(new_n1293), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1303), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1297), .B1(new_n1302), .B2(new_n1287), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  XOR2_X1   g1142(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1343));
  AOI21_X1  g1143(.A(new_n1294), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1344), .B2(new_n1331), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT127), .B1(new_n1346), .B2(new_n1330), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1304), .B1(new_n1344), .B2(new_n1337), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1343), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1332), .A2(new_n1349), .ZN(new_n1350));
  AND4_X1   g1150(.A1(KEYINPUT127), .A2(new_n1330), .A3(new_n1348), .A4(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1336), .B1(new_n1347), .B2(new_n1351), .ZN(G405));
  XNOR2_X1  g1152(.A(G375), .B(G378), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1331), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1304), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  OR2_X1    g1158(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1359), .A2(new_n1341), .A3(new_n1355), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1360), .ZN(G402));
endmodule


