

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U323 ( .A(G120GAT), .B(KEYINPUT70), .Z(n291) );
  XNOR2_X1 U324 ( .A(n350), .B(n291), .ZN(n322) );
  XNOR2_X1 U325 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U326 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n511) );
  XNOR2_X1 U327 ( .A(n512), .B(n511), .ZN(n541) );
  XNOR2_X1 U328 ( .A(G1GAT), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U329 ( .A(n292), .B(G155GAT), .ZN(n431) );
  XOR2_X1 U330 ( .A(G29GAT), .B(G134GAT), .Z(n413) );
  XOR2_X1 U331 ( .A(n431), .B(n413), .Z(n294) );
  NAND2_X1 U332 ( .A1(G225GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U334 ( .A(n295), .B(KEYINPUT1), .Z(n299) );
  XOR2_X1 U335 ( .A(G120GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n368) );
  XNOR2_X1 U338 ( .A(n368), .B(KEYINPUT5), .ZN(n298) );
  XNOR2_X1 U339 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U340 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n301) );
  XNOR2_X1 U341 ( .A(G148GAT), .B(G85GAT), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U343 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U344 ( .A(KEYINPUT85), .B(G162GAT), .Z(n305) );
  XNOR2_X1 U345 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U346 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U347 ( .A(G141GAT), .B(n306), .ZN(n390) );
  XOR2_X1 U348 ( .A(KEYINPUT88), .B(G57GAT), .Z(n308) );
  XNOR2_X1 U349 ( .A(KEYINPUT87), .B(KEYINPUT4), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U351 ( .A(n390), .B(n309), .Z(n310) );
  XNOR2_X1 U352 ( .A(n311), .B(n310), .ZN(n400) );
  XNOR2_X1 U353 ( .A(KEYINPUT90), .B(n400), .ZN(n543) );
  XOR2_X1 U354 ( .A(KEYINPUT68), .B(G92GAT), .Z(n313) );
  XNOR2_X1 U355 ( .A(G99GAT), .B(G85GAT), .ZN(n312) );
  XNOR2_X1 U356 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U357 ( .A(G106GAT), .B(n314), .Z(n424) );
  XOR2_X1 U358 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n316) );
  XNOR2_X1 U359 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U361 ( .A(n424), .B(n317), .ZN(n325) );
  XOR2_X1 U362 ( .A(G204GAT), .B(G148GAT), .Z(n382) );
  XOR2_X1 U363 ( .A(KEYINPUT13), .B(G57GAT), .Z(n319) );
  XNOR2_X1 U364 ( .A(G71GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n430) );
  XOR2_X1 U366 ( .A(n382), .B(n430), .Z(n321) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U369 ( .A(G176GAT), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U370 ( .A(n325), .B(n324), .ZN(n471) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n326) );
  XNOR2_X1 U372 ( .A(n326), .B(KEYINPUT7), .ZN(n404) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U374 ( .A(n404), .B(n439), .Z(n328) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U377 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n330) );
  XNOR2_X1 U378 ( .A(KEYINPUT29), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U380 ( .A(n332), .B(n331), .Z(n340) );
  XOR2_X1 U381 ( .A(G113GAT), .B(G50GAT), .Z(n334) );
  XNOR2_X1 U382 ( .A(G29GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U384 ( .A(G1GAT), .B(G141GAT), .Z(n336) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(G197GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n340), .B(n339), .ZN(n567) );
  NAND2_X1 U389 ( .A1(n471), .A2(n567), .ZN(n341) );
  XNOR2_X1 U390 ( .A(n341), .B(KEYINPUT71), .ZN(n456) );
  XOR2_X1 U391 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n343) );
  XNOR2_X1 U392 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U394 ( .A(G197GAT), .B(n344), .Z(n389) );
  XOR2_X1 U395 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n346) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n364) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G190GAT), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n347), .B(KEYINPUT76), .ZN(n412) );
  XNOR2_X1 U400 ( .A(n364), .B(n412), .ZN(n358) );
  XOR2_X1 U401 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n349) );
  XNOR2_X1 U402 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U404 ( .A(G8GAT), .B(G183GAT), .Z(n438) );
  XOR2_X1 U405 ( .A(n438), .B(n350), .Z(n352) );
  XNOR2_X1 U406 ( .A(G218GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U408 ( .A(n354), .B(n353), .Z(n356) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n389), .B(n359), .ZN(n540) );
  INV_X1 U413 ( .A(n540), .ZN(n491) );
  XOR2_X1 U414 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n361) );
  XNOR2_X1 U415 ( .A(G134GAT), .B(G190GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n375) );
  XOR2_X1 U417 ( .A(G99GAT), .B(G43GAT), .Z(n363) );
  NAND2_X1 U418 ( .A1(G227GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U420 ( .A(n365), .B(n364), .Z(n373) );
  XOR2_X1 U421 ( .A(KEYINPUT20), .B(G71GAT), .Z(n367) );
  XNOR2_X1 U422 ( .A(G15GAT), .B(G176GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n368), .B(G183GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n369), .B(G127GAT), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n479) );
  INV_X1 U429 ( .A(n479), .ZN(n549) );
  NAND2_X1 U430 ( .A1(n491), .A2(n549), .ZN(n392) );
  XOR2_X1 U431 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n377) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(KEYINPUT82), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U434 ( .A(G78GAT), .B(G155GAT), .Z(n379) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n387) );
  XOR2_X1 U438 ( .A(G50GAT), .B(G218GAT), .Z(n414) );
  XOR2_X1 U439 ( .A(KEYINPUT86), .B(n382), .Z(n384) );
  NAND2_X1 U440 ( .A1(G228GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n414), .B(n385), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n546) );
  NAND2_X1 U446 ( .A1(n392), .A2(n546), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT25), .ZN(n394) );
  XNOR2_X1 U448 ( .A(KEYINPUT95), .B(n394), .ZN(n398) );
  NOR2_X1 U449 ( .A1(n546), .A2(n549), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n395), .B(KEYINPUT26), .ZN(n565) );
  XOR2_X1 U451 ( .A(KEYINPUT27), .B(n540), .Z(n401) );
  NAND2_X1 U452 ( .A1(n565), .A2(n401), .ZN(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT94), .B(n396), .ZN(n397) );
  NAND2_X1 U454 ( .A1(n398), .A2(n397), .ZN(n399) );
  NAND2_X1 U455 ( .A1(n400), .A2(n399), .ZN(n403) );
  INV_X1 U456 ( .A(n543), .ZN(n489) );
  NAND2_X1 U457 ( .A1(n489), .A2(n401), .ZN(n527) );
  XOR2_X1 U458 ( .A(KEYINPUT28), .B(n546), .Z(n495) );
  NOR2_X1 U459 ( .A1(n527), .A2(n495), .ZN(n513) );
  NAND2_X1 U460 ( .A1(n513), .A2(n479), .ZN(n402) );
  NAND2_X1 U461 ( .A1(n403), .A2(n402), .ZN(n453) );
  NAND2_X1 U462 ( .A1(n404), .A2(KEYINPUT66), .ZN(n408) );
  INV_X1 U463 ( .A(n404), .ZN(n406) );
  INV_X1 U464 ( .A(KEYINPUT66), .ZN(n405) );
  NAND2_X1 U465 ( .A1(n406), .A2(n405), .ZN(n407) );
  NAND2_X1 U466 ( .A1(n408), .A2(n407), .ZN(n410) );
  AND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U472 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n418) );
  XNOR2_X1 U473 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n417) );
  XOR2_X1 U474 ( .A(n418), .B(n417), .Z(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n426) );
  XOR2_X1 U476 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n422) );
  XNOR2_X1 U477 ( .A(G162GAT), .B(KEYINPUT73), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n521) );
  XOR2_X1 U481 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n428) );
  NAND2_X1 U482 ( .A1(G231GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U484 ( .A(n429), .B(KEYINPUT12), .Z(n433) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n435) );
  XNOR2_X1 U488 ( .A(G211GAT), .B(G64GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n504) );
  INV_X1 U493 ( .A(n504), .ZN(n574) );
  NAND2_X1 U494 ( .A1(n521), .A2(n574), .ZN(n442) );
  XOR2_X1 U495 ( .A(KEYINPUT16), .B(n442), .Z(n443) );
  AND2_X1 U496 ( .A1(n453), .A2(n443), .ZN(n473) );
  NAND2_X1 U497 ( .A1(n456), .A2(n473), .ZN(n451) );
  NOR2_X1 U498 ( .A1(n543), .A2(n451), .ZN(n444) );
  XOR2_X1 U499 ( .A(KEYINPUT34), .B(n444), .Z(n445) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(n445), .ZN(G1324GAT) );
  NOR2_X1 U501 ( .A1(n540), .A2(n451), .ZN(n446) );
  XOR2_X1 U502 ( .A(G8GAT), .B(n446), .Z(G1325GAT) );
  NOR2_X1 U503 ( .A1(n451), .A2(n479), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n448) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(G1326GAT) );
  INV_X1 U508 ( .A(n495), .ZN(n482) );
  NOR2_X1 U509 ( .A1(n482), .A2(n451), .ZN(n452) );
  XOR2_X1 U510 ( .A(G22GAT), .B(n452), .Z(G1327GAT) );
  XNOR2_X1 U511 ( .A(n521), .B(KEYINPUT36), .ZN(n582) );
  NAND2_X1 U512 ( .A1(n504), .A2(n453), .ZN(n454) );
  NOR2_X1 U513 ( .A1(n582), .A2(n454), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n455), .Z(n486) );
  NAND2_X1 U515 ( .A1(n456), .A2(n486), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT38), .ZN(n458) );
  XNOR2_X1 U517 ( .A(KEYINPUT98), .B(n458), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n543), .A2(n466), .ZN(n460) );
  XNOR2_X1 U519 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  NOR2_X1 U521 ( .A1(n540), .A2(n466), .ZN(n462) );
  XNOR2_X1 U522 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(G1329GAT) );
  NOR2_X1 U524 ( .A1(n479), .A2(n466), .ZN(n464) );
  XNOR2_X1 U525 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U527 ( .A(G43GAT), .B(n465), .Z(G1330GAT) );
  NOR2_X1 U528 ( .A1(n482), .A2(n466), .ZN(n468) );
  XNOR2_X1 U529 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(G1331GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n470) );
  XNOR2_X1 U532 ( .A(G57GAT), .B(KEYINPUT103), .ZN(n469) );
  XNOR2_X1 U533 ( .A(n470), .B(n469), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT41), .B(n471), .ZN(n533) );
  XNOR2_X1 U535 ( .A(KEYINPUT102), .B(n533), .ZN(n552) );
  INV_X1 U536 ( .A(n552), .ZN(n472) );
  NOR2_X1 U537 ( .A1(n567), .A2(n472), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n473), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n543), .A2(n481), .ZN(n474) );
  XOR2_X1 U540 ( .A(n475), .B(n474), .Z(G1332GAT) );
  NOR2_X1 U541 ( .A1(n540), .A2(n481), .ZN(n477) );
  XNOR2_X1 U542 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n476) );
  XNOR2_X1 U543 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U544 ( .A(G64GAT), .B(n478), .ZN(G1333GAT) );
  NOR2_X1 U545 ( .A1(n479), .A2(n481), .ZN(n480) );
  XOR2_X1 U546 ( .A(G71GAT), .B(n480), .Z(G1334GAT) );
  NOR2_X1 U547 ( .A1(n482), .A2(n481), .ZN(n484) );
  XNOR2_X1 U548 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U550 ( .A(G78GAT), .B(n485), .Z(G1335GAT) );
  NAND2_X1 U551 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U552 ( .A(KEYINPUT108), .B(n488), .Z(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n489), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n491), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U557 ( .A(G99GAT), .B(KEYINPUT109), .Z(n494) );
  NAND2_X1 U558 ( .A1(n549), .A2(n496), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1338GAT) );
  NAND2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT44), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G106GAT), .B(n498), .ZN(G1339GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT110), .B(n504), .Z(n557) );
  NAND2_X1 U564 ( .A1(n533), .A2(n567), .ZN(n500) );
  XOR2_X1 U565 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U567 ( .A1(n521), .A2(n501), .ZN(n502) );
  NOR2_X1 U568 ( .A1(n557), .A2(n502), .ZN(n503) );
  XOR2_X1 U569 ( .A(KEYINPUT47), .B(n503), .Z(n510) );
  NOR2_X1 U570 ( .A1(n504), .A2(n582), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT45), .ZN(n506) );
  NAND2_X1 U572 ( .A1(n506), .A2(n471), .ZN(n507) );
  NOR2_X1 U573 ( .A1(n567), .A2(n507), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT112), .B(n508), .ZN(n509) );
  NOR2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n512) );
  NAND2_X1 U576 ( .A1(n549), .A2(n513), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n541), .A2(n514), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(n567), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(G120GAT), .B(KEYINPUT49), .Z(n517) );
  NAND2_X1 U581 ( .A1(n522), .A2(n552), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n519) );
  NAND2_X1 U584 ( .A1(n522), .A2(n557), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G127GAT), .B(n520), .ZN(G1342GAT) );
  XOR2_X1 U587 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  INV_X1 U588 ( .A(n521), .ZN(n560) );
  NAND2_X1 U589 ( .A1(n522), .A2(n560), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  XNOR2_X1 U591 ( .A(G141GAT), .B(KEYINPUT114), .ZN(n529) );
  INV_X1 U592 ( .A(n541), .ZN(n525) );
  NAND2_X1 U593 ( .A1(n525), .A2(n565), .ZN(n526) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n567), .A2(n537), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(G1344GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n531) );
  XNOR2_X1 U598 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(n532), .Z(n535) );
  NAND2_X1 U601 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U603 ( .A1(n574), .A2(n537), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U605 ( .A(G162GAT), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U606 ( .A1(n537), .A2(n560), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1347GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT54), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(KEYINPUT65), .ZN(n566) );
  NAND2_X1 U612 ( .A1(n566), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT55), .ZN(n548) );
  AND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n561), .A2(n567), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT57), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G183GAT), .B(n559), .ZN(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n581) );
  INV_X1 U631 ( .A(n581), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  OR2_X1 U638 ( .A1(n581), .A2(n471), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

