//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT73), .B(G902), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n190), .A2(G953), .A3(new_n187), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT21), .B(G898), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G214), .B1(G237), .B2(G902), .ZN(new_n196));
  OAI21_X1  g010(.A(G210), .B1(G237), .B2(G902), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT82), .A3(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(new_n198), .A3(KEYINPUT82), .A4(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G101), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT83), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n200), .A2(new_n213), .A3(new_n202), .A4(new_n204), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n207), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT68), .A2(G116), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT68), .A2(G116), .ZN(new_n218));
  OAI21_X1  g032(.A(G119), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n220), .A2(KEYINPUT67), .A3(G119), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT67), .B1(new_n220), .B2(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n225), .ZN(new_n227));
  INV_X1    g041(.A(new_n225), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n228), .A2(new_n219), .A3(new_n222), .A4(new_n221), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT69), .A3(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n216), .A2(KEYINPUT88), .A3(new_n226), .A4(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n226), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n205), .A2(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n232), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(G110), .B(G122), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n201), .B2(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n198), .A2(KEYINPUT84), .A3(G104), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n202), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n214), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n214), .A2(new_n245), .A3(KEYINPUT86), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G116), .ZN(new_n252));
  OAI211_X1 g066(.A(G113), .B(new_n252), .C1(new_n223), .C2(new_n250), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n248), .A2(new_n229), .A3(new_n249), .A4(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n231), .A2(new_n238), .A3(new_n240), .A4(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n231), .A2(new_n238), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n239), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n239), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT0), .A4(G128), .ZN(new_n267));
  XNOR2_X1  g081(.A(G143), .B(G146), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT90), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(G143), .B2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n265), .A2(G146), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n263), .A2(G143), .ZN(new_n277));
  OAI22_X1  g091(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n264), .A2(new_n266), .A3(new_n273), .A4(G128), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n270), .A2(new_n282), .A3(G125), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n272), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n188), .A2(G224), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n262), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n214), .A2(new_n245), .A3(KEYINPUT86), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT86), .B1(new_n214), .B2(new_n245), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n229), .A4(new_n253), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n253), .A2(new_n229), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n246), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n239), .B(KEYINPUT8), .Z(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n272), .A2(new_n300), .A3(new_n281), .A4(new_n283), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n285), .A2(KEYINPUT7), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n301), .B(new_n302), .Z(new_n303));
  AND3_X1   g117(.A1(new_n299), .A2(new_n303), .A3(new_n255), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n197), .B1(new_n288), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n286), .B1(new_n260), .B2(new_n261), .ZN(new_n307));
  INV_X1    g121(.A(new_n197), .ZN(new_n308));
  NOR4_X1   g122(.A1(new_n307), .A2(G902), .A3(new_n308), .A4(new_n304), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n195), .B(new_n196), .C1(new_n306), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G475), .ZN(new_n311));
  XNOR2_X1  g125(.A(G113), .B(G122), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n201), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n279), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(G125), .A2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(G146), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n188), .A3(G214), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n265), .ZN(new_n322));
  NOR2_X1   g136(.A1(G237), .A2(G953), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G143), .A3(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT18), .A2(G131), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND4_X1   g141(.A1(G143), .A2(new_n320), .A3(new_n188), .A4(G214), .ZN(new_n328));
  AOI21_X1  g142(.A(G143), .B1(new_n323), .B2(G214), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT93), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n331), .A3(new_n324), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT94), .A4(new_n326), .ZN(new_n336));
  AOI211_X1 g150(.A(new_n319), .B(new_n327), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n318), .A2(KEYINPUT16), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n279), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G146), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n316), .B2(new_n317), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n263), .B1(new_n343), .B2(new_n339), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT64), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n325), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n322), .A2(new_n350), .A3(new_n324), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n325), .A2(KEYINPUT17), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT95), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n325), .A2(new_n358), .A3(KEYINPUT17), .A4(new_n351), .ZN(new_n359));
  AND4_X1   g173(.A1(new_n345), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n314), .B1(new_n337), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n335), .A2(new_n336), .ZN(new_n362));
  INV_X1    g176(.A(new_n319), .ZN(new_n363));
  INV_X1    g177(.A(new_n327), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n345), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n313), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n311), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n337), .A2(new_n314), .A3(new_n360), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n318), .B(KEYINPUT19), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n263), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n341), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n352), .A2(new_n354), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n338), .A2(KEYINPUT79), .A3(G146), .A4(new_n340), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n313), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n311), .B(new_n369), .C1(new_n371), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n378), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n314), .B1(new_n337), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT96), .B1(new_n382), .B2(new_n367), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n380), .B1(KEYINPUT20), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n371), .B2(new_n379), .ZN(new_n386));
  AOI21_X1  g200(.A(G475), .B1(new_n382), .B2(new_n367), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n369), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n370), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G122), .B1(new_n217), .B2(new_n218), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n220), .A2(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n198), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT97), .B1(new_n265), .B2(G128), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT97), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n275), .A3(G143), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n397), .A2(new_n399), .B1(G128), .B2(new_n265), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n399), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n403), .B2(G134), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n265), .A2(G128), .ZN(new_n405));
  AND4_X1   g219(.A1(KEYINPUT13), .A2(new_n401), .A3(G134), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n396), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT14), .B(G122), .C1(new_n217), .C2(new_n218), .ZN(new_n408));
  OAI211_X1 g222(.A(G107), .B(new_n408), .C1(new_n393), .C2(KEYINPUT14), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n400), .A2(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(G134), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n395), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT9), .B(G234), .ZN(new_n414));
  INV_X1    g228(.A(G217), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(G953), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n407), .A2(new_n412), .A3(new_n416), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n190), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n421), .C1(KEYINPUT15), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI211_X1 g238(.A(KEYINPUT15), .B(new_n422), .C1(new_n420), .C2(new_n421), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n390), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n310), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G137), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT80), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n275), .A2(G119), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n251), .A2(G128), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT74), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n251), .A2(G128), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n275), .A2(G119), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT74), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT24), .B(G110), .Z(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT75), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n439), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n251), .B2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT23), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT23), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n436), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT77), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n450), .A3(new_n453), .A4(new_n436), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(G110), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n341), .A2(new_n344), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n445), .A2(new_n455), .A3(KEYINPUT78), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n318), .A2(new_n263), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n451), .A2(G110), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n440), .B1(new_n435), .B2(new_n439), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n375), .A2(new_n377), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n432), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n431), .B(new_n467), .C1(new_n459), .C2(new_n460), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n421), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT25), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n415), .B1(new_n421), .B2(G234), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT25), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n421), .C1(new_n469), .C2(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n469), .A2(new_n470), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n473), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n482));
  INV_X1    g296(.A(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(G134), .ZN(new_n484));
  INV_X1    g298(.A(G134), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT65), .A3(G137), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT11), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n485), .B2(G137), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(KEYINPUT11), .A3(G134), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(new_n350), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n485), .B2(G137), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n485), .A2(G137), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(KEYINPUT66), .A3(G134), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n275), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n280), .B(new_n498), .C1(new_n499), .C2(new_n268), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n498), .B1(new_n278), .B2(new_n280), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n491), .B(new_n497), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n270), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n489), .A2(new_n490), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n346), .B1(new_n506), .B2(new_n487), .ZN(new_n507));
  INV_X1    g321(.A(new_n491), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n233), .A2(new_n503), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n280), .B1(new_n499), .B2(new_n268), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n491), .A3(new_n497), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n280), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n516), .A2(G128), .B1(new_n264), .B2(new_n266), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT70), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n500), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n491), .A2(new_n497), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n485), .A2(KEYINPUT65), .A3(G137), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT65), .B1(new_n485), .B2(G137), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n524), .B2(new_n505), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n491), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n519), .A2(new_n521), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n514), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  INV_X1    g342(.A(new_n233), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n510), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n323), .A2(G210), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(G101), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n233), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n270), .B1(new_n525), .B2(new_n491), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n512), .A2(new_n491), .A3(new_n497), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n527), .A2(KEYINPUT28), .A3(new_n233), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n537), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n503), .A2(new_n509), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n549), .A3(new_n544), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n510), .A2(new_n547), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT29), .A3(new_n535), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n421), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G472), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n511), .B1(new_n503), .B2(new_n509), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT30), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n529), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n538), .A3(new_n535), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n545), .A2(new_n536), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT31), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n530), .A2(new_n563), .A3(new_n535), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n561), .A2(new_n562), .A3(new_n564), .A4(KEYINPUT71), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n556), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  AOI211_X1 g386(.A(KEYINPUT32), .B(new_n572), .C1(new_n567), .C2(new_n568), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n555), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n516), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G128), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n268), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n515), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n576), .B1(new_n582), .B2(new_n246), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n504), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n519), .A2(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n248), .A2(new_n249), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n587), .A2(new_n526), .ZN(new_n588));
  XNOR2_X1  g402(.A(G110), .B(G140), .ZN(new_n589));
  INV_X1    g403(.A(G227), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G953), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n589), .B(new_n591), .Z(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n291), .A2(new_n512), .B1(new_n246), .B2(new_n582), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT12), .A3(new_n526), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT12), .B1(new_n594), .B2(new_n526), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n526), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT87), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n587), .A2(new_n601), .A3(new_n526), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n592), .B1(new_n603), .B2(new_n588), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n575), .B(new_n421), .C1(new_n598), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n575), .A2(new_n369), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n595), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n588), .B1(new_n608), .B2(new_n596), .ZN(new_n609));
  INV_X1    g423(.A(new_n592), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n602), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n601), .B1(new_n587), .B2(new_n526), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n611), .B(G469), .C1(new_n614), .C2(new_n593), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G221), .B1(new_n414), .B2(G902), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT81), .Z(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n428), .A2(new_n481), .A3(new_n574), .A4(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(new_n213), .Z(G3));
  AOI21_X1  g436(.A(new_n190), .B1(new_n567), .B2(new_n568), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n572), .B1(new_n567), .B2(new_n568), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n480), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n620), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  INV_X1    g443(.A(new_n370), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT20), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n388), .A2(new_n386), .B1(new_n387), .B2(new_n369), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n407), .A2(new_n412), .A3(new_n416), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n416), .B1(new_n407), .B2(new_n412), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT33), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n418), .A2(new_n637), .A3(new_n419), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n422), .B1(new_n639), .B2(new_n421), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n420), .A2(new_n422), .A3(new_n421), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT99), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n190), .B1(new_n636), .B2(new_n638), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n644), .B(new_n641), .C1(new_n645), .C2(new_n422), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n310), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  XOR2_X1   g466(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n380), .B(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n426), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n630), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n310), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n629), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n625), .A2(new_n626), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n461), .A2(new_n468), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n432), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n478), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n476), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n662), .B1(new_n476), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n428), .A2(new_n620), .A3(new_n661), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G110), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  OAI21_X1  g488(.A(new_n196), .B1(new_n306), .B2(new_n309), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n189), .B1(new_n191), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n676), .A2(new_n574), .A3(new_n620), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  NAND2_X1  g495(.A1(new_n549), .A2(new_n538), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n535), .B1(new_n510), .B2(new_n547), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n535), .A2(new_n530), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n684), .B2(G902), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n571), .B2(new_n573), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n476), .A2(new_n666), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n196), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n390), .A2(new_n690), .A3(new_n426), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n306), .A2(new_n309), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(KEYINPUT38), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT38), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n306), .A2(new_n309), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n689), .A2(new_n691), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n696), .A3(KEYINPUT103), .A4(new_n691), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n678), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n620), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT40), .Z(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(new_n678), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n633), .A2(new_n647), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n676), .A2(new_n574), .A3(new_n620), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND2_X1  g523(.A1(new_n603), .A2(new_n588), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n610), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n597), .A2(new_n595), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n588), .A3(new_n592), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n421), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n619), .A3(new_n605), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n649), .A2(new_n481), .A3(new_n574), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n657), .A2(new_n481), .A3(new_n574), .A4(new_n717), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT104), .B(G116), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G18));
  NOR2_X1   g537(.A1(new_n427), .A2(new_n194), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n676), .A2(new_n574), .A3(new_n717), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  AOI21_X1  g540(.A(new_n563), .B1(new_n530), .B2(new_n535), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n520), .B1(new_n518), .B2(new_n500), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT30), .B1(new_n728), .B2(new_n541), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n233), .B1(new_n729), .B2(new_n514), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n510), .A4(new_n536), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT71), .B1(new_n732), .B2(new_n562), .ZN(new_n733));
  INV_X1    g547(.A(new_n568), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n421), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G472), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n550), .A2(KEYINPUT105), .A3(new_n551), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT105), .B1(new_n550), .B2(new_n551), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n535), .ZN(new_n739));
  INV_X1    g553(.A(new_n732), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n570), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n736), .A2(new_n481), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n310), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n633), .A2(new_n655), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n745), .A4(new_n717), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  OAI211_X1 g561(.A(new_n688), .B(new_n741), .C1(new_n623), .C2(new_n624), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n633), .A2(new_n647), .A3(new_n706), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n675), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n717), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  XNOR2_X1  g567(.A(new_n626), .B(new_n556), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n480), .B1(new_n754), .B2(new_n555), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n258), .A2(new_n239), .A3(new_n256), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n259), .B2(new_n257), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n369), .B(new_n305), .C1(new_n760), .C2(new_n286), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n308), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n288), .A2(new_n197), .A3(new_n305), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n196), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n749), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n755), .A2(new_n620), .A3(new_n758), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n574), .A3(new_n481), .A4(new_n620), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n756), .A3(new_n757), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NOR3_X1   g584(.A1(new_n764), .A2(new_n656), .A3(new_n678), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n755), .A2(new_n620), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n614), .A2(new_n593), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n592), .B1(new_n712), .B2(new_n588), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n611), .B(KEYINPUT45), .C1(new_n614), .C2(new_n593), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(G469), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT107), .A4(G469), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n606), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n605), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n785), .B(new_n606), .C1(new_n781), .C2(new_n782), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n618), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT43), .B1(new_n390), .B2(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n647), .A2(new_n390), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n688), .C1(new_n626), .C2(new_n625), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n788), .A2(new_n701), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n764), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n795), .B(new_n796), .C1(new_n793), .C2(new_n792), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT109), .B(G137), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n787), .B2(new_n618), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT47), .B(new_n619), .C1(new_n784), .C2(new_n786), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n754), .A2(new_n555), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n480), .A3(new_n804), .A4(new_n765), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  OR2_X1    g620(.A1(G952), .A2(G953), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n716), .A2(new_n605), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n808), .A2(new_n764), .A3(new_n480), .A4(new_n618), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n687), .A3(new_n189), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n811));
  INV_X1    g625(.A(new_n647), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n809), .A2(new_n687), .A3(new_n813), .A4(new_n189), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n390), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n791), .A2(new_n189), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n717), .A3(new_n796), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(new_n748), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n742), .ZN(new_n819));
  INV_X1    g633(.A(new_n696), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n690), .A3(new_n717), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(KEYINPUT117), .A3(new_n690), .A4(new_n717), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n815), .B(new_n818), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n716), .A2(new_n618), .A3(new_n605), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n801), .A2(new_n802), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n823), .A2(new_n824), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n833), .A2(new_n796), .B1(new_n834), .B2(new_n826), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n828), .B(new_n831), .C1(new_n819), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n831), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n796), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n826), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n819), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n840), .B2(new_n827), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n829), .A2(new_n830), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n811), .A2(new_n633), .A3(new_n647), .A4(new_n814), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n816), .A2(new_n751), .A3(new_n717), .A4(new_n742), .ZN(new_n844));
  AND4_X1   g658(.A1(G952), .A2(new_n843), .A3(new_n188), .A4(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n836), .A2(new_n841), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n648), .A2(KEYINPUT110), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n390), .A2(new_n655), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n633), .A2(new_n647), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n627), .A2(new_n743), .A3(new_n851), .A4(new_n620), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n621), .A2(new_n671), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n750), .A2(new_n620), .A3(new_n796), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT111), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n748), .A2(new_n764), .A3(new_n749), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(KEYINPUT111), .A3(new_n620), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n616), .A2(new_n619), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n754), .B2(new_n555), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n654), .A2(new_n426), .A3(new_n706), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n669), .A2(new_n764), .A3(new_n370), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n853), .A2(new_n859), .A3(new_n772), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n746), .A2(new_n718), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n725), .A2(new_n721), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n769), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n691), .B(new_n706), .C1(new_n306), .C2(new_n309), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n688), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n620), .A3(new_n872), .A4(new_n686), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n680), .A2(new_n708), .A3(new_n752), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n861), .B(new_n676), .C1(new_n679), .C2(new_n707), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT112), .A3(new_n752), .A4(new_n873), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n869), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT111), .B1(new_n857), .B2(new_n620), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n736), .A2(new_n707), .A3(new_n688), .A4(new_n741), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n888), .A2(new_n855), .A3(new_n860), .A4(new_n764), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n772), .B(new_n864), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n621), .A2(new_n671), .A3(new_n852), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n868), .B1(new_n865), .B2(KEYINPUT116), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n874), .A2(new_n879), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n767), .B(new_n758), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n718), .A2(new_n725), .A3(new_n746), .A4(new_n721), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n892), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n896), .B2(new_n897), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT113), .B1(new_n907), .B2(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n869), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n886), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n869), .B(new_n883), .C1(new_n880), .C2(new_n881), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n876), .A2(new_n878), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n869), .A4(new_n883), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n908), .A2(new_n911), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n846), .B(new_n902), .C1(new_n901), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n755), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n817), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n807), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n480), .A2(new_n618), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n926), .A2(new_n196), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  OR4_X1    g743(.A1(new_n686), .A2(new_n929), .A3(new_n696), .A4(new_n790), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  NOR2_X1   g745(.A1(new_n262), .A2(new_n287), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n307), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT55), .Z(new_n934));
  AOI211_X1 g748(.A(new_n421), .B(new_n197), .C1(new_n885), .C2(new_n899), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(KEYINPUT56), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n188), .A2(G952), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n885), .A2(new_n899), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n190), .A3(new_n308), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT56), .ZN(new_n941));
  INV_X1    g755(.A(new_n934), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n936), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n936), .A2(new_n943), .A3(new_n946), .A4(new_n938), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G51));
  XNOR2_X1  g762(.A(new_n606), .B(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT57), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(KEYINPUT57), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n939), .A2(KEYINPUT54), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n901), .B1(new_n885), .B2(new_n899), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n714), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n900), .A2(new_n421), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n781), .A3(new_n782), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n937), .B1(new_n955), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n956), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n382), .A2(new_n367), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n956), .A2(KEYINPUT58), .A3(G475), .A4(new_n960), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n962), .A2(new_n938), .A3(new_n963), .ZN(G60));
  OAI21_X1  g778(.A(new_n902), .B1(new_n919), .B2(new_n901), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT59), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n639), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n952), .A2(new_n953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n639), .A2(new_n968), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n969), .A2(new_n937), .A3(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n939), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n477), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n939), .A2(new_n665), .A3(new_n976), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n938), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT61), .B1(new_n980), .B2(KEYINPUT123), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G66));
  NOR2_X1   g797(.A1(new_n904), .A2(new_n891), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n188), .B1(new_n192), .B2(G224), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n760), .B1(G898), .B2(new_n188), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  AOI21_X1  g805(.A(new_n188), .B1(new_n590), .B2(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n877), .A2(new_n752), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT125), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n704), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n805), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n851), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n921), .A2(new_n702), .A3(new_n764), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n797), .A2(new_n188), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n528), .B(new_n372), .Z(new_n1005));
  NOR4_X1   g819(.A1(new_n921), .A2(new_n690), .A3(new_n692), .A4(new_n744), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n788), .A3(new_n701), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n797), .A2(new_n805), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n769), .A2(new_n772), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  NAND4_X1  g824(.A1(new_n1008), .A2(new_n188), .A3(new_n995), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1005), .A2(new_n992), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n1004), .A2(new_n1005), .B1(new_n1011), .B2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(new_n908), .A2(new_n911), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n913), .A2(new_n918), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n530), .A2(new_n536), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n531), .A2(new_n535), .ZN(new_n1020));
  AND4_X1   g834(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1008), .A2(new_n984), .A3(new_n995), .A4(new_n1010), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n1022), .B2(new_n1018), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n797), .A2(new_n984), .A3(new_n1002), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(new_n997), .A3(new_n805), .A4(new_n998), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1020), .B1(new_n1025), .B2(new_n1018), .ZN(new_n1026));
  NOR4_X1   g840(.A1(new_n1021), .A2(new_n937), .A3(new_n1023), .A4(new_n1026), .ZN(G57));
endmodule


