//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n190), .A3(G125), .ZN(new_n196));
  AOI211_X1 g010(.A(new_n188), .B(new_n189), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n188), .A2(new_n189), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT75), .A2(G146), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT89), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n196), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT75), .A3(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G237), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G214), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(G237), .A2(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(G143), .A3(G214), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT17), .A3(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n218), .A3(new_n213), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n201), .A2(new_n206), .A3(new_n215), .A4(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(G113), .B(G122), .Z(new_n222));
  XOR2_X1   g036(.A(KEYINPUT88), .B(G104), .Z(new_n223));
  XOR2_X1   g037(.A(new_n222), .B(new_n223), .Z(new_n224));
  NAND3_X1  g038(.A1(new_n214), .A2(KEYINPUT18), .A3(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n211), .A2(new_n213), .A3(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n191), .A2(new_n193), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n228), .A2(new_n189), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n189), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n225), .B(new_n227), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n221), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n221), .A2(KEYINPUT90), .A3(new_n224), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n202), .A2(new_n189), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n228), .B(KEYINPUT19), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(new_n189), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n216), .A2(new_n219), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n224), .B1(new_n241), .B2(new_n231), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n245));
  NOR2_X1   g059(.A1(G475), .A2(G902), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT91), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n236), .A2(KEYINPUT91), .A3(new_n243), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n251), .B2(KEYINPUT20), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n221), .A2(new_n231), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n236), .B1(new_n224), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G475), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n187), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT91), .B1(new_n236), .B2(new_n243), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n248), .B(new_n242), .C1(new_n234), .C2(new_n235), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n262), .B2(new_n246), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT92), .B(new_n257), .C1(new_n263), .C2(new_n247), .ZN(new_n264));
  INV_X1    g078(.A(G478), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT15), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  INV_X1    g081(.A(G116), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n268), .A2(KEYINPUT14), .A3(G122), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT14), .ZN(new_n270));
  XNOR2_X1  g084(.A(G116), .B(G122), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n267), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n210), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n274), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT95), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n276), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n274), .A2(new_n283), .ZN(new_n286));
  OAI21_X1  g100(.A(G134), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT93), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(KEYINPUT94), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n278), .A2(KEYINPUT94), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n271), .A2(new_n267), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n273), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT73), .B(G217), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G953), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n282), .A2(new_n293), .A3(new_n297), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n266), .B1(new_n302), .B2(G902), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n301), .B(new_n255), .C1(KEYINPUT15), .C2(new_n265), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n259), .A2(new_n264), .A3(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n208), .A2(G952), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT21), .B(G898), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n316), .B(KEYINPUT83), .Z(new_n317));
  OR2_X1    g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G104), .ZN(new_n324));
  INV_X1    g138(.A(G104), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n267), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(G107), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n322), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n325), .A2(KEYINPUT3), .A3(G107), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n327), .B2(KEYINPUT3), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(G104), .ZN(new_n333));
  AOI21_X1  g147(.A(G101), .B1(new_n333), .B2(G107), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT79), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n331), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n323), .A2(G104), .ZN(new_n338));
  AOI21_X1  g152(.A(G107), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n338), .A3(G107), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n322), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n330), .B1(new_n335), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n341), .B2(new_n344), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n333), .B2(G107), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n334), .A3(KEYINPUT79), .A4(new_n336), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n329), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT80), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n354));
  INV_X1    g168(.A(G119), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G116), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(G116), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n268), .A2(G119), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(G113), .B(new_n356), .C1(new_n359), .C2(new_n354), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G113), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT2), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G113), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G116), .B(G119), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n360), .B2(new_n361), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n348), .A2(new_n353), .A3(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(G110), .B(G122), .Z(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n336), .B(new_n343), .C1(new_n339), .C2(new_n340), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(G101), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n335), .B2(new_n345), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n375), .A3(G101), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n359), .A2(KEYINPUT67), .A3(new_n364), .A4(new_n366), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT67), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n367), .B1(new_n368), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n372), .A2(new_n374), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n189), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n210), .A2(G146), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(G128), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT65), .B1(new_n189), .B2(G143), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n210), .A3(G146), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n390), .A2(new_n392), .B1(G143), .B2(new_n189), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n275), .B1(new_n386), .B2(KEYINPUT1), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n192), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n210), .B2(G146), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n189), .A2(KEYINPUT65), .A3(G143), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n386), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT0), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n275), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n399), .A3(new_n275), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n386), .A2(new_n387), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n398), .A2(new_n404), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n395), .B1(new_n406), .B2(new_n192), .ZN(new_n407));
  INV_X1    g221(.A(G224), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n408), .B2(G953), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n360), .A2(new_n369), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n352), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n373), .B(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n346), .B2(new_n371), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n410), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n385), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n321), .B1(new_n418), .B2(new_n255), .ZN(new_n419));
  AOI211_X1 g233(.A(KEYINPUT87), .B(G902), .C1(new_n385), .C2(new_n417), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n352), .A2(KEYINPUT80), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n347), .B(new_n329), .C1(new_n349), .C2(new_n351), .ZN(new_n423));
  INV_X1    g237(.A(new_n371), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n384), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n373), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(new_n373), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n408), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n407), .B(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n320), .B1(new_n421), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n319), .C1(new_n419), .C2(new_n420), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n318), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n208), .A2(G227), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n277), .B2(G137), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n277), .A2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT66), .A2(G131), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n446), .A2(new_n448), .A3(new_n451), .A4(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT10), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n422), .A2(new_n423), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n379), .A2(new_n406), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n378), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n389), .B1(new_n405), .B2(new_n394), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n329), .B(new_n462), .C1(new_n349), .C2(new_n351), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(KEYINPUT10), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n455), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n457), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n348), .A2(new_n353), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n455), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n349), .A2(new_n351), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n330), .A3(new_n461), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n470), .A2(new_n471), .B1(new_n378), .B2(new_n459), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n444), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n456), .B1(new_n469), .B2(new_n330), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT12), .B(new_n455), .C1(new_n476), .C2(new_n463), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT81), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n352), .B2(new_n456), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT81), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT12), .A4(new_n455), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n455), .B1(new_n476), .B2(new_n463), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n478), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n473), .A2(new_n444), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n474), .A2(new_n475), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n468), .B1(new_n467), .B2(new_n472), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n475), .B(new_n443), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n440), .B(new_n255), .C1(new_n487), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n440), .A2(new_n255), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n478), .A2(new_n481), .A3(new_n484), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n473), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n443), .B(KEYINPUT77), .Z(new_n496));
  AND2_X1   g310(.A1(new_n473), .A2(new_n444), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(new_n496), .B1(new_n465), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n493), .B1(new_n498), .B2(G469), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n439), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n406), .A2(new_n455), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n447), .A2(G134), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n218), .B1(new_n503), .B2(new_n449), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(new_n218), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n456), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n502), .B1(new_n501), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n383), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT68), .B1(new_n380), .B2(new_n382), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n406), .A2(new_n455), .B1(new_n506), .B2(new_n456), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n212), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n510), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n510), .A2(KEYINPUT31), .A3(new_n516), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n521), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n514), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n501), .A2(new_n531), .A3(new_n507), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n501), .A2(new_n507), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT68), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n511), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n501), .A2(new_n507), .B1(new_n382), .B2(new_n380), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n528), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NOR2_X1   g358(.A1(G472), .A2(G902), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT72), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n526), .B2(new_n527), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT32), .B1(new_n549), .B2(new_n546), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n521), .B1(new_n534), .B2(new_n540), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n510), .A2(new_n516), .A3(new_n521), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n535), .A2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n516), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT28), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n557), .A2(new_n534), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n521), .A2(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n255), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n548), .A2(new_n550), .B1(G472), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT23), .B1(new_n275), .B2(G119), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT74), .B1(new_n275), .B2(G119), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT76), .B(G110), .Z(new_n567));
  XNOR2_X1  g381(.A(G119), .B(G128), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT24), .B(G110), .Z(new_n569));
  OAI22_X1  g383(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n237), .A2(new_n229), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(G110), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n568), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n205), .A3(new_n203), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n208), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n575), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n563), .B1(new_n583), .B2(G902), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n581), .A2(KEYINPUT25), .A3(new_n255), .A4(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n295), .B1(G234), .B2(new_n255), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n583), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n587), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n562), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n307), .A2(new_n437), .A3(new_n500), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND2_X1  g409(.A1(new_n492), .A2(new_n499), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n549), .A2(new_n546), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n528), .B2(new_n542), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(KEYINPUT96), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n598), .B2(KEYINPUT96), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n596), .A2(new_n438), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n592), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n301), .A2(new_n265), .A3(new_n255), .ZN(new_n605));
  NAND2_X1  g419(.A1(G478), .A2(G902), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n301), .B(KEYINPUT33), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n265), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n259), .B2(new_n264), .ZN(new_n609));
  INV_X1    g423(.A(new_n316), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n610), .B(new_n315), .C1(new_n434), .C2(new_n436), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n603), .A2(new_n604), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND2_X1  g429(.A1(new_n251), .A2(KEYINPUT20), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n262), .A2(new_n245), .A3(new_n246), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n618), .A2(new_n257), .A3(new_n305), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n604), .A2(new_n603), .A3(new_n611), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n267), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NOR2_X1   g437(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n576), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n590), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n588), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n603), .A2(new_n307), .A3(new_n437), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  OR2_X1    g446(.A1(new_n312), .A2(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n310), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n618), .A2(new_n257), .A3(new_n305), .A4(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n610), .B1(new_n434), .B2(new_n436), .ZN(new_n637));
  INV_X1    g451(.A(new_n629), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n562), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(new_n500), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  NAND2_X1  g455(.A1(new_n259), .A2(new_n264), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n305), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n643), .A2(new_n610), .A3(new_n629), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n434), .A2(new_n436), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n548), .A2(new_n550), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n510), .A2(new_n516), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(new_n521), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n556), .A2(new_n529), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(G902), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n600), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n649), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  AOI211_X1 g471(.A(KEYINPUT100), .B(new_n655), .C1(new_n548), .C2(new_n550), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n634), .B(KEYINPUT39), .Z(new_n661));
  AOI211_X1 g475(.A(new_n439), .B(new_n661), .C1(new_n492), .C2(new_n499), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n644), .A2(new_n645), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n646), .A2(new_n660), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  INV_X1    g480(.A(new_n608), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n642), .A2(new_n667), .A3(new_n637), .A4(new_n634), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n500), .A2(new_n639), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n609), .A2(new_n672), .A3(new_n637), .A4(new_n634), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT103), .B(G146), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G48));
  OAI21_X1  g490(.A(new_n443), .B1(new_n488), .B2(new_n489), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT82), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n497), .A2(new_n494), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n490), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n440), .A3(new_n255), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n440), .B1(new_n680), .B2(new_n255), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n681), .A2(new_n682), .A3(new_n439), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n611), .A3(new_n609), .A4(new_n593), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND4_X1  g500(.A1(new_n683), .A2(new_n611), .A3(new_n593), .A4(new_n619), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT104), .B(G116), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G18));
  NOR3_X1   g503(.A1(new_n562), .A2(new_n315), .A3(new_n638), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n307), .A2(new_n683), .A3(new_n637), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  AOI21_X1  g506(.A(new_n306), .B1(new_n259), .B2(new_n264), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n637), .B1(new_n693), .B2(KEYINPUT107), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n695), .B(new_n306), .C1(new_n259), .C2(new_n264), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n681), .A2(new_n682), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n588), .A2(KEYINPUT106), .A3(new_n591), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  INV_X1    g513(.A(new_n587), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n584), .B2(new_n585), .ZN(new_n701));
  INV_X1    g515(.A(new_n591), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n528), .B1(new_n529), .B2(new_n558), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n546), .B(KEYINPUT105), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n549), .B2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n705), .A2(new_n315), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n697), .A2(new_n438), .A3(new_n711), .ZN(new_n712));
  OR3_X1    g526(.A1(new_n694), .A2(new_n696), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n638), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n697), .A2(new_n438), .A3(new_n637), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n609), .A2(new_n634), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n192), .ZN(G27));
  XNOR2_X1  g533(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n647), .B2(new_n610), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n434), .A2(new_n722), .A3(new_n436), .A4(new_n316), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n493), .B(KEYINPUT108), .Z(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n498), .B2(G469), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n439), .B1(new_n492), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n593), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n720), .B1(new_n728), .B2(new_n717), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n721), .A2(new_n723), .A3(new_n727), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n562), .A2(new_n705), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n609), .A2(new_n634), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NOR2_X1   g550(.A1(new_n728), .A2(new_n635), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT111), .B(G134), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G36));
  NAND2_X1  g553(.A1(new_n498), .A2(KEYINPUT45), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  INV_X1    g555(.A(new_n496), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n494), .B2(new_n473), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n486), .A2(new_n489), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n724), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n724), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n492), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n438), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n661), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n721), .A2(new_n723), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n259), .A2(new_n667), .A3(new_n264), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n259), .A2(new_n264), .A3(new_n667), .A4(new_n760), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n602), .B(new_n638), .C1(new_n758), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n755), .B1(KEYINPUT44), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n762), .B2(KEYINPUT44), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n752), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n438), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n634), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n608), .B(new_n773), .C1(new_n259), .C2(new_n264), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n562), .A2(new_n754), .A3(new_n592), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND2_X1  g591(.A1(new_n680), .A2(new_n255), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G469), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n438), .A3(new_n492), .ZN(new_n780));
  AOI21_X1  g594(.A(G902), .B1(new_n385), .B2(new_n417), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n321), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n319), .B1(new_n782), .B2(new_n435), .ZN(new_n783));
  INV_X1    g597(.A(new_n436), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n316), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n715), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n780), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n635), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n787), .A2(new_n774), .B1(new_n671), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n643), .A2(new_n695), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n629), .B2(new_n773), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n628), .A2(KEYINPUT115), .A3(new_n588), .A4(new_n634), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n657), .B2(new_n658), .ZN(new_n795));
  INV_X1    g609(.A(new_n727), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n790), .A2(new_n797), .A3(new_n637), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n674), .A2(new_n789), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n674), .A2(new_n789), .A3(new_n799), .A4(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT116), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n727), .B(new_n794), .C1(new_n658), .C2(new_n657), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n694), .A2(new_n696), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT52), .B(new_n640), .C1(new_n716), .C2(new_n717), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n809), .B2(new_n674), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n802), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n594), .A2(new_n687), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n500), .A2(new_n437), .A3(new_n604), .A4(new_n602), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n667), .B1(new_n259), .B2(new_n264), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n307), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n630), .A2(new_n684), .A3(new_n691), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n727), .A2(new_n715), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n305), .A2(new_n773), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n618), .A2(new_n819), .A3(new_n257), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n618), .A2(new_n819), .A3(KEYINPUT114), .A4(new_n257), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n717), .A2(new_n818), .B1(new_n824), .B2(new_n670), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n754), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n816), .A2(new_n817), .A3(new_n713), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n737), .B1(new_n729), .B2(new_n734), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n811), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n800), .A2(new_n801), .B1(new_n809), .B2(new_n674), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n642), .A2(new_n608), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n642), .B2(new_n305), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n594), .B(new_n687), .C1(new_n834), .C2(new_n813), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n630), .A2(new_n684), .A3(new_n691), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n828), .A3(new_n713), .A4(new_n826), .ZN(new_n838));
  XOR2_X1   g652(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n839));
  NOR3_X1   g653(.A1(new_n832), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT54), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n811), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n839), .B1(new_n832), .B2(new_n838), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n310), .B1(new_n758), .B2(new_n761), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n754), .A3(new_n683), .A4(new_n715), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n659), .A2(new_n310), .A3(new_n592), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n642), .A2(new_n667), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n683), .A3(new_n754), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n697), .A2(new_n439), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n770), .A2(new_n771), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n705), .A2(new_n710), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n849), .A2(new_n857), .A3(new_n754), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n648), .A2(new_n316), .A3(new_n780), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n857), .A3(new_n849), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(KEYINPUT50), .A3(new_n857), .A4(new_n849), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n866), .A2(KEYINPUT118), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n866), .B2(KEYINPUT118), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n562), .A2(new_n705), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n849), .A2(new_n754), .A3(new_n683), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT48), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n849), .A2(new_n637), .A3(new_n683), .A4(new_n857), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n851), .A2(new_n609), .A3(new_n683), .A4(new_n754), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n308), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n868), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n848), .A2(new_n876), .B1(G952), .B2(G953), .ZN(new_n877));
  OR4_X1    g691(.A1(new_n317), .A2(new_n659), .A3(new_n439), .A4(new_n705), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n697), .B(KEYINPUT49), .Z(new_n879));
  OR4_X1    g693(.A1(new_n648), .A2(new_n878), .A3(new_n756), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(new_n880), .ZN(G75));
  NOR2_X1   g695(.A1(new_n208), .A2(G952), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n694), .A2(new_n696), .A3(new_n712), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n835), .A2(new_n836), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n826), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n803), .A2(KEYINPUT116), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n809), .A2(new_n805), .A3(new_n674), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n802), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n839), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n802), .A2(new_n803), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n830), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(G210), .B(G902), .C1(new_n889), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n428), .A2(new_n430), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n432), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n882), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n844), .A2(new_n846), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT120), .A3(G210), .A4(G902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n900), .A2(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n724), .B(KEYINPUT57), .Z(new_n908));
  NOR3_X1   g722(.A1(new_n889), .A2(new_n892), .A3(KEYINPUT54), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n680), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n889), .A2(new_n892), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n913), .A2(new_n255), .A3(new_n746), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n882), .B1(new_n912), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  OAI211_X1 g730(.A(G902), .B(new_n916), .C1(new_n889), .C2(new_n892), .ZN(new_n917));
  INV_X1    g731(.A(new_n262), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n882), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n918), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT121), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G60));
  XOR2_X1   g738(.A(new_n606), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n607), .B1(new_n848), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n607), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n909), .B2(new_n910), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n920), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n625), .B(new_n934), .C1(new_n889), .C2(new_n892), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n882), .B1(KEYINPUT122), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n844), .B2(new_n846), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n935), .B(new_n937), .C1(new_n938), .C2(new_n589), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT123), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n583), .B1(new_n913), .B2(new_n933), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n941), .A3(new_n935), .A4(new_n937), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(G66));
  NOR2_X1   g760(.A1(new_n314), .A2(new_n408), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n208), .ZN(new_n948));
  INV_X1    g762(.A(new_n884), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n208), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n896), .B1(G898), .B2(new_n208), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(G69));
  AOI21_X1  g766(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n515), .B(new_n502), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n238), .ZN(new_n955));
  NAND2_X1  g769(.A1(G900), .A2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n694), .A2(new_n696), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n753), .A2(new_n957), .A3(new_n870), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n674), .A2(new_n789), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n829), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n767), .A2(new_n776), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n955), .B(new_n956), .C1(new_n961), .C2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  INV_X1    g778(.A(new_n665), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n959), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n665), .A2(KEYINPUT62), .A3(new_n674), .A4(new_n789), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n307), .A2(new_n814), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n754), .A2(new_n969), .A3(new_n593), .A4(new_n662), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n772), .B2(new_n775), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n767), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n955), .B1(new_n973), .B2(new_n208), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n953), .B1(new_n963), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n953), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n973), .A2(new_n208), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n976), .B(new_n962), .C1(new_n977), .C2(new_n955), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(G72));
  XNOR2_X1  g793(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n980));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n973), .B2(new_n949), .ZN(new_n983));
  INV_X1    g797(.A(new_n652), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n961), .B2(new_n949), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n882), .B1(new_n986), .B2(new_n553), .ZN(new_n987));
  INV_X1    g801(.A(new_n553), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n652), .A2(new_n988), .A3(new_n982), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT126), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n831), .B2(new_n840), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n985), .A2(new_n987), .A3(new_n991), .ZN(G57));
endmodule


