

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(KEYINPUT97), .ZN(n792) );
  NOR2_X1 U551 ( .A1(n784), .A2(n773), .ZN(n515) );
  AND2_X1 U552 ( .A1(n765), .A2(n764), .ZN(n516) );
  INV_X1 U553 ( .A(KEYINPUT30), .ZN(n714) );
  XNOR2_X1 U554 ( .A(n714), .B(KEYINPUT93), .ZN(n715) );
  XNOR2_X1 U555 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U556 ( .A1(n706), .A2(n705), .ZN(n749) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n706) );
  NOR2_X1 U558 ( .A1(G651), .A2(n643), .ZN(n638) );
  XOR2_X1 U559 ( .A(n517), .B(KEYINPUT17), .Z(n870) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  NAND2_X1 U561 ( .A1(n870), .A2(G137), .ZN(n520) );
  INV_X1 U562 ( .A(G2105), .ZN(n521) );
  AND2_X1 U563 ( .A1(n521), .A2(G2104), .ZN(n871) );
  NAND2_X1 U564 ( .A1(G101), .A2(n871), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U566 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n866) );
  NAND2_X1 U568 ( .A1(G113), .A2(n866), .ZN(n523) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n521), .ZN(n867) );
  NAND2_X1 U570 ( .A1(G125), .A2(n867), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U572 ( .A1(n525), .A2(n524), .ZN(G160) );
  NAND2_X1 U573 ( .A1(G138), .A2(n870), .ZN(n532) );
  NAND2_X1 U574 ( .A1(n866), .A2(G114), .ZN(n526) );
  XOR2_X1 U575 ( .A(n526), .B(KEYINPUT82), .Z(n530) );
  NAND2_X1 U576 ( .A1(G102), .A2(n871), .ZN(n528) );
  NAND2_X1 U577 ( .A1(G126), .A2(n867), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(G164) );
  INV_X1 U581 ( .A(G651), .ZN(n536) );
  NOR2_X1 U582 ( .A1(G543), .A2(n536), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n533), .Z(n642) );
  NAND2_X1 U584 ( .A1(G64), .A2(n642), .ZN(n535) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  NAND2_X1 U586 ( .A1(G52), .A2(n638), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n629) );
  NAND2_X1 U589 ( .A1(G90), .A2(n629), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n643), .A2(n536), .ZN(n630) );
  NAND2_X1 U591 ( .A1(G77), .A2(n630), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(G171) );
  NAND2_X1 U595 ( .A1(G135), .A2(n870), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n542), .B(KEYINPUT74), .ZN(n549) );
  NAND2_X1 U597 ( .A1(G111), .A2(n866), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G99), .A2(n871), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n867), .A2(G123), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT18), .B(n545), .Z(n546) );
  NOR2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n993) );
  XNOR2_X1 U604 ( .A(G2096), .B(n993), .ZN(n550) );
  OR2_X1 U605 ( .A1(G2100), .A2(n550), .ZN(G156) );
  NAND2_X1 U606 ( .A1(G65), .A2(n642), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G53), .A2(n638), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G91), .A2(n629), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G78), .A2(n630), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n729) );
  INV_X1 U613 ( .A(n729), .ZN(G299) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  NAND2_X1 U615 ( .A1(G88), .A2(n629), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G75), .A2(n630), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G62), .A2(n642), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G50), .A2(n638), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G166) );
  NAND2_X1 U622 ( .A1(n629), .A2(G89), .ZN(n563) );
  XNOR2_X1 U623 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G76), .A2(n630), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U627 ( .A1(G63), .A2(n642), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G51), .A2(n638), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT71), .ZN(G286) );
  NAND2_X1 U635 ( .A1(G94), .A2(G452), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT65), .ZN(G173) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U638 ( .A(n575), .B(KEYINPUT66), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT10), .B(n576), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n813) );
  NAND2_X1 U641 ( .A1(n813), .A2(G567), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U643 ( .A1(G81), .A2(n629), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT68), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U646 ( .A1(G68), .A2(n630), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n582), .Z(n586) );
  NAND2_X1 U649 ( .A1(G56), .A2(n642), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT67), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n584), .B(KEYINPUT14), .ZN(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n638), .A2(G43), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n971) );
  INV_X1 U655 ( .A(G860), .ZN(n604) );
  OR2_X1 U656 ( .A1(n971), .A2(n604), .ZN(G153) );
  INV_X1 U657 ( .A(G171), .ZN(G301) );
  NAND2_X1 U658 ( .A1(G79), .A2(n630), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G54), .A2(n638), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G92), .A2(n629), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G66), .A2(n642), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT69), .B(n593), .Z(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT15), .B(n596), .ZN(n976) );
  NOR2_X1 U667 ( .A1(G868), .A2(n976), .ZN(n598) );
  INV_X1 U668 ( .A(G868), .ZN(n601) );
  NOR2_X1 U669 ( .A1(n601), .A2(G301), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U671 ( .A(KEYINPUT70), .B(n599), .ZN(G284) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n600), .B(KEYINPUT72), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n601), .A2(G286), .ZN(n602) );
  NOR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n604), .A2(G559), .ZN(n605) );
  INV_X1 U677 ( .A(n976), .ZN(n885) );
  NAND2_X1 U678 ( .A1(n605), .A2(n885), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n971), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n885), .A2(G868), .ZN(n607) );
  NOR2_X1 U682 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT73), .B(n610), .Z(G282) );
  NAND2_X1 U685 ( .A1(n885), .A2(G559), .ZN(n655) );
  XNOR2_X1 U686 ( .A(n971), .B(n655), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n611), .A2(G860), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G55), .A2(n638), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT76), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G93), .A2(n629), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT75), .B(n613), .Z(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G80), .A2(n630), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G67), .A2(n642), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n649) );
  XNOR2_X1 U697 ( .A(n620), .B(n649), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G73), .A2(n630), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G61), .A2(n642), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G48), .A2(n638), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n629), .A2(G86), .ZN(n624) );
  XOR2_X1 U704 ( .A(KEYINPUT78), .B(n624), .Z(n625) );
  NOR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(G305) );
  NAND2_X1 U707 ( .A1(G85), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G72), .A2(n630), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G60), .A2(n642), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G47), .A2(n638), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT64), .B(n637), .Z(G290) );
  NAND2_X1 U715 ( .A1(G49), .A2(n638), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G87), .A2(n643), .ZN(n644) );
  XOR2_X1 U720 ( .A(KEYINPUT77), .B(n644), .Z(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(G288) );
  NOR2_X1 U722 ( .A1(G868), .A2(n649), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n647), .B(KEYINPUT79), .ZN(n658) );
  XOR2_X1 U724 ( .A(G305), .B(n971), .Z(n648) );
  XOR2_X1 U725 ( .A(n649), .B(n648), .Z(n650) );
  XOR2_X1 U726 ( .A(n650), .B(KEYINPUT19), .Z(n652) );
  XNOR2_X1 U727 ( .A(G290), .B(G166), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(G299), .ZN(n884) );
  XNOR2_X1 U731 ( .A(n884), .B(n655), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n664) );
  NAND2_X1 U741 ( .A1(G132), .A2(G82), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(KEYINPUT80), .ZN(n666) );
  NOR2_X1 U744 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(G96), .A2(n667), .ZN(n819) );
  NAND2_X1 U746 ( .A1(G2106), .A2(n819), .ZN(n671) );
  NAND2_X1 U747 ( .A1(G120), .A2(G69), .ZN(n668) );
  NOR2_X1 U748 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(G108), .A2(n669), .ZN(n820) );
  NAND2_X1 U750 ( .A1(G567), .A2(n820), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n842) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U753 ( .A1(n842), .A2(n672), .ZN(n816) );
  NAND2_X1 U754 ( .A1(n816), .A2(G36), .ZN(G176) );
  INV_X1 U755 ( .A(G166), .ZN(G303) );
  AND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n705) );
  INV_X1 U757 ( .A(n705), .ZN(n674) );
  NOR2_X1 U758 ( .A1(n706), .A2(n674), .ZN(n808) );
  NAND2_X1 U759 ( .A1(G140), .A2(n870), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G104), .A2(n871), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U762 ( .A(KEYINPUT34), .B(n677), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G116), .A2(n866), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G128), .A2(n867), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U766 ( .A(KEYINPUT83), .B(n680), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT35), .B(n681), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT36), .B(n684), .ZN(n853) );
  XNOR2_X1 U770 ( .A(KEYINPUT37), .B(G2067), .ZN(n796) );
  NOR2_X1 U771 ( .A1(n853), .A2(n796), .ZN(n996) );
  NAND2_X1 U772 ( .A1(n808), .A2(n996), .ZN(n803) );
  NAND2_X1 U773 ( .A1(n871), .A2(G95), .ZN(n685) );
  XNOR2_X1 U774 ( .A(n685), .B(KEYINPUT84), .ZN(n687) );
  NAND2_X1 U775 ( .A1(G131), .A2(n870), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U777 ( .A(KEYINPUT85), .B(n688), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G107), .A2(n866), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G119), .A2(n867), .ZN(n689) );
  AND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n863) );
  AND2_X1 U782 ( .A1(n863), .A2(G1991), .ZN(n704) );
  NAND2_X1 U783 ( .A1(G141), .A2(n870), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n693), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U785 ( .A1(G105), .A2(n871), .ZN(n694) );
  XOR2_X1 U786 ( .A(KEYINPUT87), .B(n694), .Z(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT38), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G117), .A2(n866), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n867), .A2(G129), .ZN(n698) );
  XOR2_X1 U791 ( .A(KEYINPUT86), .B(n698), .Z(n699) );
  NOR2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n852) );
  AND2_X1 U794 ( .A1(n852), .A2(G1996), .ZN(n703) );
  OR2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n989) );
  NAND2_X1 U796 ( .A1(n989), .A2(n808), .ZN(n797) );
  NAND2_X1 U797 ( .A1(n803), .A2(n797), .ZN(n791) );
  NAND2_X1 U798 ( .A1(G8), .A2(n749), .ZN(n784) );
  NOR2_X1 U799 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NAND2_X1 U800 ( .A1(KEYINPUT33), .A2(n959), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n784), .A2(n707), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n708), .B(KEYINPUT95), .ZN(n710) );
  XOR2_X1 U803 ( .A(KEYINPUT96), .B(G1981), .Z(n709) );
  XNOR2_X1 U804 ( .A(G305), .B(n709), .ZN(n979) );
  NAND2_X1 U805 ( .A1(n710), .A2(n979), .ZN(n777) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n749), .ZN(n763) );
  NOR2_X1 U807 ( .A1(n784), .A2(G1966), .ZN(n711) );
  XNOR2_X1 U808 ( .A(n711), .B(KEYINPUT90), .ZN(n766) );
  NOR2_X1 U809 ( .A1(n763), .A2(n766), .ZN(n712) );
  XNOR2_X1 U810 ( .A(KEYINPUT92), .B(n712), .ZN(n713) );
  NAND2_X1 U811 ( .A1(n713), .A2(G8), .ZN(n716) );
  NOR2_X1 U812 ( .A1(G168), .A2(n717), .ZN(n721) );
  XNOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NOR2_X1 U814 ( .A1(n749), .A2(n912), .ZN(n719) );
  INV_X1 U815 ( .A(n749), .ZN(n734) );
  INV_X1 U816 ( .A(G1961), .ZN(n928) );
  NOR2_X1 U817 ( .A1(n734), .A2(n928), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U819 ( .A1(G171), .A2(n723), .ZN(n720) );
  NOR2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n722), .Z(n764) );
  NAND2_X1 U822 ( .A1(G171), .A2(n723), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n734), .A2(G2072), .ZN(n724) );
  XNOR2_X1 U824 ( .A(n724), .B(KEYINPUT27), .ZN(n726) );
  XNOR2_X1 U825 ( .A(G1956), .B(KEYINPUT91), .ZN(n938) );
  NOR2_X1 U826 ( .A1(n938), .A2(n734), .ZN(n725) );
  NOR2_X1 U827 ( .A1(n726), .A2(n725), .ZN(n728) );
  NOR2_X1 U828 ( .A1(n729), .A2(n728), .ZN(n727) );
  XOR2_X1 U829 ( .A(n727), .B(KEYINPUT28), .Z(n745) );
  NAND2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n743) );
  AND2_X1 U831 ( .A1(n734), .A2(G1996), .ZN(n730) );
  XOR2_X1 U832 ( .A(n730), .B(KEYINPUT26), .Z(n732) );
  NAND2_X1 U833 ( .A1(n749), .A2(G1341), .ZN(n731) );
  NAND2_X1 U834 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U835 ( .A1(n971), .A2(n733), .ZN(n738) );
  NAND2_X1 U836 ( .A1(G1348), .A2(n749), .ZN(n736) );
  NAND2_X1 U837 ( .A1(G2067), .A2(n734), .ZN(n735) );
  NAND2_X1 U838 ( .A1(n736), .A2(n735), .ZN(n739) );
  NOR2_X1 U839 ( .A1(n976), .A2(n739), .ZN(n737) );
  OR2_X1 U840 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U841 ( .A1(n976), .A2(n739), .ZN(n740) );
  NAND2_X1 U842 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U844 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U845 ( .A(KEYINPUT29), .B(n746), .Z(n747) );
  NAND2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n765) );
  INV_X1 U847 ( .A(G8), .ZN(n755) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n784), .ZN(n751) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U850 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U851 ( .A(n752), .B(KEYINPUT94), .ZN(n753) );
  NAND2_X1 U852 ( .A1(n753), .A2(G303), .ZN(n754) );
  OR2_X1 U853 ( .A1(n755), .A2(n754), .ZN(n757) );
  AND2_X1 U854 ( .A1(n765), .A2(n757), .ZN(n756) );
  NAND2_X1 U855 ( .A1(n764), .A2(n756), .ZN(n761) );
  INV_X1 U856 ( .A(n757), .ZN(n759) );
  AND2_X1 U857 ( .A1(G286), .A2(G8), .ZN(n758) );
  OR2_X1 U858 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U859 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U860 ( .A(n762), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G8), .A2(n763), .ZN(n768) );
  NOR2_X1 U862 ( .A1(n516), .A2(n766), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n783) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U866 ( .A1(n959), .A2(n771), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n783), .A2(n772), .ZN(n774) );
  NAND2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n960) );
  INV_X1 U869 ( .A(n960), .ZN(n773) );
  AND2_X1 U870 ( .A1(n774), .A2(n515), .ZN(n775) );
  NOR2_X1 U871 ( .A1(KEYINPUT33), .A2(n775), .ZN(n776) );
  NOR2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U874 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  NOR2_X1 U875 ( .A1(n784), .A2(n779), .ZN(n780) );
  XNOR2_X1 U876 ( .A(n780), .B(KEYINPUT89), .ZN(n787) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U878 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n793) );
  XNOR2_X1 U884 ( .A(n793), .B(n792), .ZN(n795) );
  XNOR2_X1 U885 ( .A(G290), .B(G1986), .ZN(n964) );
  NAND2_X1 U886 ( .A1(n964), .A2(n808), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n811) );
  AND2_X1 U888 ( .A1(n853), .A2(n796), .ZN(n990) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n852), .ZN(n1005) );
  INV_X1 U890 ( .A(n797), .ZN(n800) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n863), .ZN(n992) );
  NOR2_X1 U892 ( .A1(G290), .A2(G1986), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n992), .A2(n798), .ZN(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n1005), .A2(n801), .ZN(n802) );
  XNOR2_X1 U896 ( .A(KEYINPUT39), .B(n802), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT98), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n990), .A2(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(KEYINPUT99), .B(n807), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U907 ( .A1(G3), .A2(G1), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT101), .B(n815), .Z(n817) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT102), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  INV_X1 U913 ( .A(G132), .ZN(G219) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  INV_X1 U916 ( .A(G82), .ZN(G220) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  XOR2_X1 U919 ( .A(G1966), .B(G1981), .Z(n822) );
  XNOR2_X1 U920 ( .A(G1996), .B(G1991), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n822), .B(n821), .ZN(n832) );
  XOR2_X1 U922 ( .A(KEYINPUT108), .B(G2474), .Z(n824) );
  XNOR2_X1 U923 ( .A(G1961), .B(KEYINPUT106), .ZN(n823) );
  XNOR2_X1 U924 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U925 ( .A(G1971), .B(G1956), .Z(n826) );
  XNOR2_X1 U926 ( .A(G1986), .B(G1976), .ZN(n825) );
  XNOR2_X1 U927 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U928 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U929 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(G229) );
  XOR2_X1 U932 ( .A(KEYINPUT105), .B(G2084), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2078), .B(G2072), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(G2100), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(G227) );
  XOR2_X1 U942 ( .A(KEYINPUT104), .B(n842), .Z(G319) );
  NAND2_X1 U943 ( .A1(G112), .A2(n866), .ZN(n844) );
  NAND2_X1 U944 ( .A1(G100), .A2(n871), .ZN(n843) );
  NAND2_X1 U945 ( .A1(n844), .A2(n843), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n870), .A2(G136), .ZN(n845) );
  XNOR2_X1 U947 ( .A(KEYINPUT109), .B(n845), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n867), .A2(G124), .ZN(n846) );
  XOR2_X1 U949 ( .A(KEYINPUT44), .B(n846), .Z(n847) );
  NOR2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(KEYINPUT110), .B(n849), .Z(n850) );
  NOR2_X1 U952 ( .A1(n851), .A2(n850), .ZN(G162) );
  XOR2_X1 U953 ( .A(n853), .B(n852), .Z(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(n993), .ZN(n862) );
  NAND2_X1 U955 ( .A1(G139), .A2(n870), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G103), .A2(n871), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G115), .A2(n866), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G127), .A2(n867), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(KEYINPUT47), .B(n859), .Z(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n1000) );
  XOR2_X1 U963 ( .A(n862), .B(n1000), .Z(n865) );
  XOR2_X1 U964 ( .A(G160), .B(n863), .Z(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n879) );
  NAND2_X1 U966 ( .A1(G118), .A2(n866), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G130), .A2(n867), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G142), .A2(n870), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G106), .A2(n871), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U972 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U974 ( .A(KEYINPUT48), .B(n877), .Z(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U976 ( .A(G164), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n882), .B(G162), .ZN(n883) );
  NOR2_X1 U979 ( .A1(G37), .A2(n883), .ZN(G395) );
  XOR2_X1 U980 ( .A(n884), .B(G286), .Z(n887) );
  XNOR2_X1 U981 ( .A(G171), .B(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G37), .A2(n888), .ZN(G397) );
  NOR2_X1 U984 ( .A1(G229), .A2(G227), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n889), .B(KEYINPUT49), .ZN(n902) );
  XOR2_X1 U986 ( .A(G2443), .B(G2427), .Z(n891) );
  XNOR2_X1 U987 ( .A(G2438), .B(G2454), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(n892), .B(G2435), .Z(n894) );
  XNOR2_X1 U990 ( .A(G1341), .B(G1348), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U992 ( .A(G2430), .B(G2446), .Z(n896) );
  XNOR2_X1 U993 ( .A(KEYINPUT100), .B(G2451), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n898), .B(n897), .Z(n899) );
  NAND2_X1 U996 ( .A1(G14), .A2(n899), .ZN(n905) );
  NAND2_X1 U997 ( .A1(n905), .A2(G319), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT111), .B(n900), .Z(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  INV_X1 U1004 ( .A(n905), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n1018) );
  XOR2_X1 U1006 ( .A(G29), .B(KEYINPUT114), .Z(n925) );
  XOR2_X1 U1007 ( .A(G2072), .B(G33), .Z(n906) );
  NAND2_X1 U1008 ( .A1(n906), .A2(G28), .ZN(n909) );
  XOR2_X1 U1009 ( .A(KEYINPUT113), .B(G1996), .Z(n907) );
  XNOR2_X1 U1010 ( .A(G32), .B(n907), .ZN(n908) );
  NOR2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n916) );
  XOR2_X1 U1012 ( .A(G2067), .B(G26), .Z(n911) );
  XOR2_X1 U1013 ( .A(G1991), .B(G25), .Z(n910) );
  NAND2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n914) );
  XOR2_X1 U1015 ( .A(G27), .B(n912), .Z(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT53), .ZN(n920) );
  XOR2_X1 U1019 ( .A(G2084), .B(G34), .Z(n918) );
  XNOR2_X1 U1020 ( .A(KEYINPUT54), .B(n918), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G35), .B(G2090), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT55), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n926), .A2(G11), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT115), .B(n927), .Z(n958) );
  XNOR2_X1 U1028 ( .A(n928), .B(G5), .ZN(n951) );
  XOR2_X1 U1029 ( .A(G1966), .B(G21), .Z(n937) );
  XOR2_X1 U1030 ( .A(G1986), .B(G24), .Z(n931) );
  XOR2_X1 U1031 ( .A(G22), .B(KEYINPUT120), .Z(n929) );
  XNOR2_X1 U1032 ( .A(n929), .B(G1971), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT121), .B(G1976), .Z(n932) );
  XNOR2_X1 U1035 ( .A(G23), .B(n932), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(n935), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n949) );
  XOR2_X1 U1039 ( .A(n938), .B(G20), .Z(n942) );
  XNOR2_X1 U1040 ( .A(G1348), .B(G4), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(n939), .B(KEYINPUT119), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(KEYINPUT59), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G19), .B(G1341), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n947), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n952), .B(KEYINPUT123), .ZN(n954) );
  XOR2_X1 U1052 ( .A(KEYINPUT61), .B(KEYINPUT122), .Z(n953) );
  XNOR2_X1 U1053 ( .A(n954), .B(n953), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(G16), .A2(n955), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(n956), .B(KEYINPUT124), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n987) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n985) );
  INV_X1 U1058 ( .A(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1060 ( .A(KEYINPUT117), .B(n962), .Z(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G166), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n965), .B(KEYINPUT118), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G1956), .B(KEYINPUT116), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(n966), .B(G299), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G301), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G1341), .B(n971), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G1348), .B(n976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT57), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(KEYINPUT125), .ZN(n1016) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n999) );
  XOR2_X1 U1082 ( .A(G160), .B(G2084), .Z(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(KEYINPUT112), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1010) );
  XOR2_X1 U1088 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n1003), .ZN(n1008) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n1006), .Z(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1011), .ZN(n1013) );
  INV_X1 U1098 ( .A(KEYINPUT55), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1018), .B(n1017), .ZN(G150) );
  INV_X1 U1103 ( .A(G150), .ZN(G311) );
endmodule

