//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n217), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n216), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G20), .A2(G77), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT15), .B(G87), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT72), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n223), .A2(G33), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n247), .B1(new_n249), .B2(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n222), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT66), .A2(G1), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(G13), .A3(G20), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT66), .A2(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT66), .A2(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n268), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n257), .B1(new_n265), .B2(new_n269), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G77), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n222), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G107), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n209), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(new_n232), .A3(G1698), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n277), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n261), .A2(new_n291), .A3(new_n262), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT67), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n268), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n277), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G244), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  AND2_X1   g0098(.A1(G1), .A2(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n260), .A3(new_n291), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n288), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(G200), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(new_n274), .A3(new_n271), .A4(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n278), .A2(G222), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G223), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n315), .B1(new_n258), .B2(new_n278), .C1(new_n279), .C2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(new_n277), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT65), .B(G226), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n296), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n305), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n324));
  INV_X1    g0124(.A(G58), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT8), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(KEYINPUT68), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n254), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n223), .A2(KEYINPUT69), .A3(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n323), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n257), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n272), .A2(G50), .A3(new_n273), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n270), .A2(new_n202), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n318), .A2(new_n337), .A3(new_n320), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n322), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n322), .A2(KEYINPUT71), .A3(new_n336), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n278), .A2(G226), .A3(new_n314), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n313), .B1(new_n347), .B2(new_n277), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n296), .A2(G238), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n331), .B2(new_n258), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n257), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT11), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n360), .A3(new_n257), .ZN(new_n361));
  INV_X1    g0161(.A(new_n273), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n208), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n359), .A2(new_n361), .B1(new_n272), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n265), .A2(new_n269), .A3(new_n208), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n355), .B(new_n368), .C1(new_n308), .C2(new_n354), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n312), .A2(new_n343), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n371), .A3(new_n366), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n364), .B2(new_n366), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n352), .B1(new_n348), .B2(new_n349), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(G169), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n337), .B2(new_n354), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n376), .B1(new_n354), .B2(G169), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n375), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n318), .B2(new_n320), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n336), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n387), .B(new_n389), .C1(new_n308), .C2(new_n321), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n336), .B2(new_n388), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n384), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n392), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n318), .A2(new_n320), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n386), .B1(G190), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n384), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n389), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n370), .A2(new_n383), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n286), .B2(new_n223), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n402), .B(G20), .C1(new_n283), .C2(new_n285), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT75), .B1(G58), .B2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(G58), .C2(G68), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n278), .B2(G20), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n208), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n407), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n415), .A2(new_n405), .A3(new_n201), .ZN(new_n416));
  INV_X1    g0216(.A(G159), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n416), .A2(new_n223), .B1(new_n417), .B2(new_n249), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n411), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n419), .A3(new_n257), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n327), .A2(new_n362), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n272), .B1(new_n270), .B2(new_n327), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n313), .B1(new_n296), .B2(G232), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n278), .A2(G226), .A3(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n278), .A2(G223), .A3(new_n314), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n282), .C2(new_n210), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n277), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G190), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n296), .A2(G232), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n428), .A3(new_n302), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n423), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n420), .A2(new_n422), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n424), .A2(new_n337), .A3(new_n428), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n305), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n437), .A2(KEYINPUT18), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n441));
  AOI21_X1  g0241(.A(G169), .B1(new_n424), .B2(new_n428), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n337), .B2(new_n429), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT18), .A4(new_n437), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n438), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n423), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n441), .A2(new_n445), .A3(new_n448), .A4(KEYINPUT77), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n436), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n400), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n284), .A2(G33), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n457));
  OAI21_X1  g0257(.A(G303), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n283), .A2(new_n285), .A3(G264), .A4(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n283), .A2(new_n285), .A3(G257), .A4(new_n314), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT83), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(KEYINPUT83), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n277), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(G274), .B1(new_n276), .B2(new_n222), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n261), .A2(G45), .A3(new_n262), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n266), .A2(new_n267), .A3(new_n290), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n277), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(G270), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT21), .A3(G169), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n465), .A2(G179), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n256), .A2(new_n222), .B1(G20), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G20), .B1(G33), .B2(G283), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n282), .A2(G97), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT85), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT85), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT20), .B(new_n481), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(new_n489), .B1(new_n270), .B2(new_n480), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n265), .A2(new_n269), .ZN(new_n491));
  INV_X1    g0291(.A(new_n257), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n268), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n491), .A2(G116), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT84), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n272), .A2(new_n496), .A3(G116), .A4(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n479), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n305), .B1(new_n465), .B2(new_n475), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n490), .A2(new_n495), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n476), .A2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n465), .A2(G190), .A3(new_n475), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(new_n497), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n499), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n278), .A2(new_n510), .A3(new_n223), .A4(G87), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n283), .A2(new_n285), .A3(new_n223), .A4(G87), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  INV_X1    g0316(.A(new_n254), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n223), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n280), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n517), .A2(G116), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n515), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n515), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n257), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n272), .A2(new_n493), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n491), .B2(G107), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n265), .A2(new_n269), .A3(KEYINPUT25), .A4(new_n280), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n525), .A2(G107), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n283), .A2(new_n285), .A3(G257), .A4(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n283), .A2(new_n285), .A3(G250), .A4(new_n314), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G294), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n277), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n472), .A2(new_n473), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n299), .A2(new_n300), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(G264), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n472), .A2(new_n301), .A3(new_n473), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n534), .A2(new_n537), .A3(new_n538), .A4(new_n308), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT88), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n534), .A2(new_n537), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT87), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n471), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT87), .ZN(new_n545));
  AOI21_X1  g0345(.A(G200), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n524), .B(new_n529), .C1(new_n541), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(G179), .A3(new_n545), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n542), .B2(new_n471), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n529), .A2(new_n524), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n535), .A2(KEYINPUT78), .A3(G257), .A4(new_n536), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(new_n536), .C1(new_n467), .C2(new_n470), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n283), .A2(new_n285), .A3(G250), .A4(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(new_n314), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n277), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n565), .A3(new_n538), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G169), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n558), .A2(new_n565), .A3(G179), .A4(new_n538), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n401), .B2(new_n403), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT6), .ZN(new_n571));
  AND2_X1   g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n280), .A2(KEYINPUT6), .A3(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G97), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n578), .A2(new_n257), .B1(new_n579), .B2(new_n270), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n272), .A2(G97), .A3(new_n493), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT79), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n248), .A2(G77), .ZN(new_n583));
  INV_X1    g0383(.A(new_n575), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(new_n571), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n583), .B1(new_n586), .B2(new_n223), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n280), .B1(new_n412), .B2(new_n413), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n257), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n270), .A2(new_n579), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(new_n581), .A3(KEYINPUT79), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n569), .B1(new_n582), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n558), .A2(new_n565), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(G190), .A3(new_n538), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n566), .A2(G200), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n581), .A3(new_n580), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n272), .A2(G87), .A3(new_n493), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n270), .A2(new_n253), .ZN(new_n599));
  NAND3_X1  g0399(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n223), .A2(new_n600), .B1(new_n573), .B2(new_n210), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT81), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n283), .A2(new_n285), .A3(new_n223), .A4(G68), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n254), .B2(new_n579), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n601), .C2(new_n602), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n257), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n598), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT80), .B1(new_n466), .B2(new_n467), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT80), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n472), .A2(new_n612), .A3(new_n301), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n283), .A2(new_n285), .A3(G238), .A4(new_n314), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(G1698), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G116), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n277), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n277), .A2(new_n211), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n467), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n614), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n614), .A2(new_n619), .A3(G190), .A4(new_n621), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n610), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n611), .A2(new_n613), .B1(new_n467), .B2(new_n620), .ZN(new_n626));
  AOI21_X1  g0426(.A(G169), .B1(new_n626), .B2(new_n619), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n614), .A2(new_n619), .A3(new_n621), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n337), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT82), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(new_n223), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n573), .A2(new_n210), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT81), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n603), .A3(new_n605), .A4(new_n607), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n257), .A2(new_n635), .B1(new_n270), .B2(new_n253), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n251), .B(KEYINPUT72), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n491), .A2(new_n637), .A3(new_n492), .A4(new_n493), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n630), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n630), .A2(new_n638), .A3(new_n599), .A4(new_n609), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n629), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n593), .A2(new_n597), .A3(new_n625), .A4(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n455), .A2(new_n509), .A3(new_n553), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n448), .A2(new_n440), .ZN(new_n644));
  INV_X1    g0444(.A(new_n307), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n383), .B1(new_n369), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n646), .B2(new_n436), .ZN(new_n647));
  INV_X1    g0447(.A(new_n399), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n341), .B2(new_n342), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n626), .A2(new_n337), .A3(new_n619), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n628), .B2(G169), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n638), .A2(new_n599), .A3(new_n609), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT82), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n636), .A2(new_n630), .A3(new_n638), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n624), .A2(new_n598), .A3(new_n599), .A4(new_n609), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT89), .B(new_n385), .C1(new_n626), .C2(new_n619), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n622), .B2(G200), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT90), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n623), .A2(KEYINPUT89), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n622), .A2(new_n658), .A3(G200), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n610), .A3(new_n624), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n641), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n589), .A2(new_n581), .A3(new_n590), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n569), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT26), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT79), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n673), .A2(new_n591), .B1(new_n567), .B2(new_n568), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n625), .A3(new_n641), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n656), .B1(G200), .B2(new_n622), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n655), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n674), .A4(new_n676), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n552), .A2(new_n499), .A3(new_n503), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n673), .A2(new_n591), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n668), .B1(G200), .B2(new_n566), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n569), .A2(new_n686), .B1(new_n687), .B2(new_n595), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n547), .A3(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n641), .A2(new_n662), .A3(new_n665), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n662), .B1(new_n641), .B2(new_n665), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n641), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n649), .B1(new_n454), .B2(new_n694), .ZN(G369));
  AND2_X1   g0495(.A1(new_n508), .A2(KEYINPUT93), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n223), .A2(G13), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n268), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n498), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n508), .B2(KEYINPUT93), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n497), .A2(new_n504), .B1(new_n477), .B2(new_n478), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT21), .B1(new_n498), .B2(new_n500), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n696), .A2(new_n705), .B1(new_n708), .B2(new_n704), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n551), .A2(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n553), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n703), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n552), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n708), .A2(new_n703), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n548), .A2(new_n549), .B1(new_n529), .B2(new_n524), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(new_n553), .B1(new_n718), .B2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  NOR2_X1   g0520(.A1(new_n632), .A2(G116), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n226), .A2(new_n289), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n220), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n676), .B1(new_n680), .B2(new_n674), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n669), .B1(new_n661), .B2(new_n666), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n706), .A2(new_n718), .A3(new_n707), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n547), .A2(new_n593), .A3(new_n597), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n655), .B1(new_n732), .B2(new_n667), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n703), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n678), .B(new_n682), .C1(new_n727), .C2(KEYINPUT26), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n703), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(KEYINPUT29), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n642), .A2(new_n509), .A3(new_n553), .A4(new_n714), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n544), .A2(new_n545), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n628), .A2(new_n558), .A3(new_n565), .ZN(new_n742));
  INV_X1    g0542(.A(new_n478), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n741), .A2(KEYINPUT30), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n594), .A2(new_n544), .A3(new_n545), .A4(new_n628), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n478), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n628), .A2(G179), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n740), .A2(new_n476), .A3(new_n748), .A4(new_n566), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n703), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n739), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n725), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n710), .A2(G330), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n697), .B(KEYINPUT95), .Z(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G45), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G1), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n760), .B(new_n711), .C1(new_n722), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n722), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n278), .A2(new_n226), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n226), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n242), .A2(new_n290), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n286), .A2(new_n226), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n221), .B2(new_n290), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n222), .B1(G20), .B2(new_n305), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n767), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n223), .A2(G179), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n210), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n223), .A2(new_n337), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n308), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n782), .A2(new_n308), .A3(G200), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n788), .A2(new_n202), .B1(new_n789), .B2(new_n280), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n223), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n784), .B(new_n790), .C1(G97), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n785), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(G190), .A3(new_n385), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n278), .B1(new_n796), .B2(new_n258), .C1(new_n325), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT32), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n782), .A2(new_n795), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n417), .ZN(new_n801));
  INV_X1    g0601(.A(new_n800), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(KEYINPUT32), .A3(G159), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n798), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n786), .A2(G190), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(KEYINPUT96), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(KEYINPUT96), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n794), .B(new_n804), .C1(new_n208), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT97), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n812), .A2(new_n789), .B1(new_n783), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n797), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G322), .B1(new_n802), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n286), .C1(new_n817), .C2(new_n796), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n788), .A2(new_n819), .B1(new_n820), .B2(new_n792), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n814), .B(new_n818), .C1(KEYINPUT98), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT33), .B(G317), .Z(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(KEYINPUT98), .B2(new_n821), .C1(new_n808), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n809), .A2(new_n810), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n811), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n781), .B1(new_n826), .B2(new_n778), .ZN(new_n827));
  INV_X1    g0627(.A(new_n777), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n710), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n765), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n275), .A2(new_n703), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n311), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n307), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n645), .A2(new_n714), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n737), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n312), .A2(new_n714), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n733), .B2(new_n736), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n838), .A2(new_n756), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n756), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n767), .B(new_n841), .C1(new_n845), .C2(KEYINPUT102), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT102), .B2(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(new_n778), .ZN(new_n848));
  INV_X1    g0648(.A(new_n808), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G283), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n797), .A2(new_n820), .B1(new_n800), .B2(new_n817), .ZN(new_n851));
  INV_X1    g0651(.A(new_n796), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n278), .B(new_n851), .C1(G116), .C2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G97), .A2(new_n793), .B1(new_n787), .B2(G303), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n789), .A2(new_n210), .ZN(new_n855));
  INV_X1    g0655(.A(new_n783), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(G107), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n850), .A2(new_n853), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n278), .B1(new_n800), .B2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n792), .A2(new_n325), .B1(new_n783), .B2(new_n202), .ZN(new_n861));
  INV_X1    g0661(.A(new_n789), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n861), .C1(G68), .C2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n815), .A2(G143), .B1(new_n852), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n865), .B2(new_n788), .C1(new_n808), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n868), .B2(KEYINPUT34), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n858), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n848), .B1(new_n872), .B2(KEYINPUT101), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(KEYINPUT101), .B2(new_n872), .ZN(new_n874));
  INV_X1    g0674(.A(new_n767), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n778), .A2(new_n775), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT100), .Z(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n258), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n874), .B(new_n879), .C1(new_n776), .C2(new_n837), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n847), .A2(new_n880), .ZN(G384));
  OR2_X1    g0681(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(G116), .A4(new_n224), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  NAND4_X1  g0685(.A1(new_n221), .A2(G77), .A3(new_n406), .A4(new_n407), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n202), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(G13), .B(new_n268), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(G330), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n382), .A2(KEYINPUT104), .ZN(new_n891));
  INV_X1    g0691(.A(new_n374), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n372), .A3(new_n703), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n369), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n375), .B(new_n895), .C1(new_n380), .C2(new_n381), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n380), .A2(new_n381), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n369), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n375), .A3(new_n703), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n755), .A3(new_n837), .ZN(new_n902));
  INV_X1    g0702(.A(new_n701), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n437), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n434), .B(new_n904), .C1(new_n423), .C2(new_n447), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n453), .B2(new_n904), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT38), .B(new_n906), .C1(new_n453), .C2(new_n904), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n905), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n434), .B(KEYINPUT17), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n904), .B1(new_n915), .B2(new_n644), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n901), .A2(new_n755), .A3(new_n837), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n455), .A2(new_n755), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n890), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  INV_X1    g0724(.A(new_n839), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n684), .B2(new_n693), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT103), .A3(new_n836), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  INV_X1    g0728(.A(new_n836), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n840), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n909), .A2(new_n910), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n901), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n891), .A2(new_n896), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n703), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n448), .A2(new_n440), .A3(new_n701), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n735), .B(new_n455), .C1(KEYINPUT29), .C2(new_n737), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n649), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n924), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n268), .B2(new_n761), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n924), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n889), .B1(new_n946), .B2(new_n947), .ZN(G367));
  NOR2_X1   g0748(.A1(new_n808), .A2(new_n820), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G283), .A2(new_n852), .B1(new_n802), .B2(G317), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n278), .B1(new_n815), .B2(G303), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n856), .A2(KEYINPUT46), .A3(G116), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n783), .B2(new_n480), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n789), .A2(new_n579), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n788), .A2(new_n817), .B1(new_n280), .B2(new_n792), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n949), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT109), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n808), .A2(new_n417), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n796), .A2(new_n202), .B1(new_n800), .B2(new_n865), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n286), .B(new_n961), .C1(G150), .C2(new_n815), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n862), .A2(G77), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n793), .A2(G68), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n787), .A2(G143), .B1(new_n856), .B2(G58), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n959), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT110), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n778), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n610), .A2(new_n714), .ZN(new_n971));
  MUX2_X1   g0771(.A(new_n692), .B(new_n641), .S(new_n971), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n777), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n779), .B1(new_n253), .B2(new_n226), .C1(new_n238), .C2(new_n772), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n767), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n763), .B(KEYINPUT108), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n668), .A2(new_n703), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n688), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n670), .A2(new_n703), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n719), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT44), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n719), .A2(new_n980), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT45), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n716), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT106), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT106), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n716), .A2(new_n985), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n717), .A2(new_n553), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n715), .B2(new_n717), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n991), .B(new_n993), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n758), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n758), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n722), .B(KEYINPUT41), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n976), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT43), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n972), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n980), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n992), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT42), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n674), .B1(new_n980), .B2(new_n718), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n703), .B1(new_n1006), .B2(KEYINPUT105), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT105), .B2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1002), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n972), .A2(new_n1001), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n716), .A2(new_n1003), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1011), .B(new_n1012), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n975), .B1(new_n1000), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT111), .ZN(G387));
  AOI21_X1  g0815(.A(new_n722), .B1(new_n994), .B2(new_n758), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n758), .B2(new_n994), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n715), .A2(new_n828), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n768), .A2(new_n721), .B1(G107), .B2(new_n226), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n235), .A2(new_n290), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n721), .ZN(new_n1021));
  AOI211_X1 g0821(.A(G45), .B(new_n1021), .C1(G68), .C2(G77), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n250), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n772), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1019), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n767), .B1(new_n1026), .B2(new_n780), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n792), .A2(new_n812), .B1(new_n783), .B2(new_n820), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n815), .A2(G317), .B1(new_n852), .B2(G303), .ZN(new_n1029));
  INV_X1    g0829(.A(G322), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n788), .C1(new_n808), .C2(new_n817), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n286), .B1(new_n800), .B2(new_n819), .C1(new_n480), .C2(new_n789), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT112), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n808), .A2(new_n327), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n783), .A2(new_n258), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n956), .B(new_n1041), .C1(G159), .C2(new_n787), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n637), .A2(new_n793), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n286), .B1(new_n802), .B2(G150), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n815), .A2(G50), .B1(new_n852), .B2(G68), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1036), .A2(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1027), .B1(new_n1047), .B2(new_n778), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n994), .A2(new_n976), .B1(new_n1018), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1017), .A2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n986), .A2(new_n989), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n995), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n996), .A2(new_n766), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n976), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1003), .A2(new_n777), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT113), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n779), .B1(new_n579), .B2(new_n226), .C1(new_n245), .C2(new_n772), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n767), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n783), .A2(new_n208), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n855), .B(new_n1060), .C1(G77), .C2(new_n793), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n286), .B1(new_n802), .B2(G143), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n250), .B2(new_n796), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n808), .C2(new_n202), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n787), .B1(new_n815), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n286), .B1(new_n800), .B2(new_n1030), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G294), .B2(new_n852), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n280), .A2(new_n789), .B1(new_n783), .B2(new_n812), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G116), .B2(new_n793), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n808), .C2(new_n813), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G317), .A2(new_n787), .B1(new_n815), .B2(G311), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1065), .A2(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1059), .B1(new_n1075), .B2(new_n778), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1057), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1053), .A2(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n843), .A2(new_n1079), .A3(new_n455), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT115), .B1(new_n756), .B2(new_n454), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1082), .A2(new_n942), .A3(new_n649), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT116), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n755), .A2(G330), .A3(new_n837), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n897), .A2(new_n900), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n901), .A2(new_n755), .A3(G330), .A4(new_n837), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n931), .A2(new_n1084), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n714), .B(new_n835), .C1(new_n693), .C2(new_n728), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n836), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n927), .A2(new_n930), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n1084), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1083), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n934), .A2(new_n936), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1086), .B1(new_n927), .B2(new_n930), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n938), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT114), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n938), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n918), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1086), .B1(new_n1092), .B2(new_n836), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1093), .A2(new_n901), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n938), .B1(new_n910), .B2(new_n917), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1088), .B1(new_n1103), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1103), .A2(new_n1112), .A3(new_n1088), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1100), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1113), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1082), .A2(new_n942), .A3(new_n649), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1097), .A2(new_n1084), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n931), .A2(new_n1089), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n722), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1116), .A2(new_n976), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n875), .B1(new_n327), .B2(new_n878), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n792), .A2(new_n258), .B1(new_n797), .B2(new_n480), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n849), .C2(G107), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n208), .A2(new_n789), .B1(new_n783), .B2(new_n210), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n286), .B1(new_n800), .B2(new_n820), .C1(new_n579), .C2(new_n796), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(G283), .C2(new_n787), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n788), .A2(new_n1133), .B1(new_n417), .B2(new_n792), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n815), .A2(G132), .B1(new_n802), .B2(G125), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  AOI21_X1  g0936(.A(new_n286), .B1(new_n852), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1134), .B(new_n1138), .C1(G50), .C2(new_n862), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT53), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n783), .B2(new_n866), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n856), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n849), .A2(G137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1129), .A2(new_n1132), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n934), .A2(new_n936), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1125), .B1(new_n848), .B2(new_n1144), .C1(new_n1145), .C2(new_n776), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1124), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1124), .A2(KEYINPUT119), .A3(new_n1146), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1123), .B1(new_n1148), .B2(new_n1149), .ZN(G378));
  OAI211_X1 g0950(.A(G330), .B(new_n920), .C1(new_n911), .C2(KEYINPUT40), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n336), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n648), .B(new_n339), .C1(new_n1152), .C2(new_n701), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n339), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n336), .B(new_n903), .C1(new_n399), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n941), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1158), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n912), .A2(G330), .A3(new_n920), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n939), .A2(new_n940), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1163), .A2(new_n1164), .B1(new_n1165), .B2(new_n933), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1162), .A2(new_n776), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n876), .A2(new_n202), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n797), .A2(new_n1133), .B1(new_n796), .B2(new_n865), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G150), .B2(new_n793), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n787), .A2(G125), .B1(new_n856), .B2(new_n1136), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n808), .C2(new_n859), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n862), .A2(G159), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1041), .B1(G58), .B2(new_n862), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n480), .B2(new_n788), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n278), .A2(G41), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n812), .B2(new_n800), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n797), .A2(new_n280), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT120), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G68), .C2(new_n793), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n253), .B2(new_n796), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1180), .B(new_n1186), .C1(G97), .C2(new_n849), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1181), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1191));
  AND4_X1   g0991(.A1(new_n1178), .A2(new_n1188), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n767), .B(new_n1169), .C1(new_n1192), .C2(new_n848), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1167), .A2(new_n1054), .B1(new_n1168), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT121), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n938), .B1(new_n931), .B2(new_n901), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1106), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT114), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1196), .A2(new_n1145), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1088), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1103), .A2(new_n1112), .A3(new_n1088), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1121), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1083), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n941), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1163), .A2(new_n933), .A3(new_n1165), .A4(new_n1164), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1195), .B1(new_n1209), .B2(new_n766), .ZN(new_n1210));
  AOI211_X1 g1010(.A(KEYINPUT121), .B(new_n722), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT122), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1203), .A2(new_n1083), .B1(new_n1207), .B2(new_n1206), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(KEYINPUT57), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1117), .B1(new_n1116), .B2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(KEYINPUT122), .B(new_n1205), .C1(new_n1218), .C2(new_n1167), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1194), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(G375));
  NAND3_X1  g1022(.A1(new_n1118), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1100), .A2(new_n999), .A3(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT123), .Z(new_n1225));
  NAND3_X1  g1025(.A1(new_n1217), .A2(KEYINPUT124), .A3(new_n976), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n767), .B1(G68), .B2(new_n877), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n849), .A2(G116), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n963), .B1(new_n788), .B2(new_n820), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G97), .B2(new_n856), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n796), .A2(new_n280), .B1(new_n800), .B2(new_n813), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n278), .B(new_n1231), .C1(G283), .C2(new_n815), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1228), .A2(new_n1043), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n849), .A2(new_n1136), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n278), .B1(new_n797), .B2(new_n865), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G150), .B2(new_n852), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n787), .A2(G132), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n793), .A2(G50), .B1(new_n862), .B2(G58), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n783), .A2(new_n417), .B1(new_n800), .B2(new_n1133), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT125), .Z(new_n1241));
  OAI21_X1  g1041(.A(new_n1233), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1227), .B1(new_n1242), .B2(new_n778), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n901), .B2(new_n776), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1216), .B2(new_n1054), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1226), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1225), .A2(new_n1247), .ZN(G381));
  NAND2_X1  g1048(.A1(new_n1123), .A2(new_n1147), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1017), .A2(new_n1049), .A3(new_n831), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G384), .A2(G390), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(G375), .A3(G381), .A4(new_n1251), .ZN(G407));
  INV_X1    g1052(.A(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n702), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1221), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1250), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G390), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT111), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1258), .B2(new_n1250), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1262), .B2(G390), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n1014), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n722), .B1(new_n1266), .B2(new_n1223), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1216), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1223), .B1(new_n1121), .B2(new_n1270), .ZN(new_n1271));
  AND4_X1   g1071(.A1(KEYINPUT126), .A2(new_n1271), .A3(new_n766), .A4(new_n1268), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1247), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G384), .B(new_n1247), .C1(new_n1269), .C2(new_n1272), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1255), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1214), .A2(new_n999), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1194), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1249), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1221), .B2(G378), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1280), .B1(new_n1284), .B2(new_n1255), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n766), .B1(new_n1218), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT121), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1209), .A2(new_n1195), .A3(new_n766), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1215), .A4(new_n1219), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G378), .A3(new_n1282), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1282), .A2(new_n1281), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1253), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1254), .A4(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1285), .A2(new_n1286), .A3(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1255), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1265), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1295), .A2(new_n1254), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1297), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1280), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1298), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1264), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(G405));
  NOR2_X1   g1111(.A1(new_n1221), .A2(new_n1249), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1292), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1298), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1298), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1265), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1264), .A3(new_n1314), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(G402));
endmodule


