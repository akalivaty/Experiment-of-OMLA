//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XOR2_X1   g036(.A(KEYINPUT3), .B(G2104), .Z(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n478), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT65), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g062(.A1(KEYINPUT65), .A2(G100), .A3(G2105), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AOI21_X1  g066(.A(new_n475), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(G126), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT66), .B(G114), .ZN(new_n495));
  OAI211_X1 g070(.A(G2104), .B(new_n494), .C1(new_n495), .C2(new_n483), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n483), .A2(G138), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n474), .A2(new_n476), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n474), .A2(KEYINPUT67), .A3(new_n476), .A4(new_n498), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n483), .A2(G138), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n497), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT68), .B(G89), .Z(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(G651), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G63), .B1(new_n510), .B2(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n531), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n510), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n515), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n518), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NOR2_X1   g114(.A1(new_n527), .A2(new_n528), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(G68), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n546));
  INV_X1    g121(.A(new_n515), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G81), .B1(G43), .B2(new_n510), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT71), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT72), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n510), .A2(G53), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n558), .B2(KEYINPUT9), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n518), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n513), .A2(new_n514), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n566), .B1(new_n571), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n564), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  OAI211_X1 g151(.A(KEYINPUT76), .B(G651), .C1(new_n514), .C2(G74), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  NAND2_X1  g153(.A1(G74), .A2(G651), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n529), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n510), .A2(G49), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n570), .C2(new_n583), .ZN(G288));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n510), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n510), .A2(new_n585), .A3(G48), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n567), .A2(G86), .A3(new_n569), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n540), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n547), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n518), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n571), .A2(G92), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT10), .Z(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n540), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g185(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g191(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g192(.A(G323), .B(new_n617), .ZN(G282));
  NOR3_X1   g193(.A1(new_n462), .A2(new_n467), .A3(G2105), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n483), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n623), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AND2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G32), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n468), .A2(G105), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  INV_X1    g257(.A(G141), .ZN(new_n683));
  INV_X1    g258(.A(new_n478), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n484), .A2(G129), .ZN(new_n686));
  NAND3_X1  g261(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT26), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n680), .B1(new_n693), .B2(new_n679), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT27), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1996), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n478), .A2(G139), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n698));
  NAND3_X1  g273(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G127), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G115), .B2(G2104), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n697), .B(new_n700), .C1(new_n703), .C2(new_n483), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n679), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n679), .B2(G33), .ZN(new_n707));
  INV_X1    g282(.A(G2072), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n629), .A2(new_n679), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT94), .Z(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NOR2_X1   g288(.A1(G171), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G5), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G28), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT30), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n719), .B2(KEYINPUT30), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n712), .A2(new_n717), .A3(new_n718), .A4(new_n724), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n709), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G164), .A2(new_n679), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G27), .B2(new_n679), .ZN(new_n728));
  INV_X1    g303(.A(G2078), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G168), .A2(new_n713), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n713), .B2(G21), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT93), .B(G1966), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n728), .A2(new_n729), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n480), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR4_X1   g318(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n696), .A2(new_n726), .A3(new_n730), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n713), .A2(G22), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT87), .Z(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G303), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n713), .A2(G6), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G305), .B2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n713), .A2(G23), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G288), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT33), .B(G1976), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n754), .A2(new_n755), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n758), .A2(new_n759), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n752), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT34), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G24), .ZN(new_n768));
  XNOR2_X1  g343(.A(G290), .B(KEYINPUT86), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1986), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n679), .A2(G25), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n478), .A2(G131), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT84), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n483), .A2(G107), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n484), .A2(G119), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n773), .B1(new_n782), .B2(new_n679), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT35), .B(G1991), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT85), .Z(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n783), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n766), .A2(new_n767), .A3(new_n772), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n713), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n551), .B2(new_n713), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n713), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n679), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n679), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT29), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n799), .B1(G2090), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n713), .A2(G4), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n607), .B2(new_n713), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1348), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n679), .A2(G26), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT28), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n478), .A2(G140), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n484), .A2(G128), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n483), .A2(G116), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n811), .B1(new_n816), .B2(G29), .ZN(new_n817));
  INV_X1    g392(.A(G2067), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n804), .A2(new_n806), .A3(new_n809), .A4(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n747), .A2(new_n790), .A3(new_n791), .A4(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n510), .A2(G55), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n515), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n518), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G860), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n607), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT38), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n549), .A2(new_n828), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT97), .Z(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n550), .B2(new_n828), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n829), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(new_n781), .B(KEYINPUT101), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n621), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n483), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n484), .A2(G130), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  AOI211_X1 g423(.A(new_n846), .B(new_n848), .C1(G142), .C2(new_n478), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n843), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n690), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n705), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n692), .B2(new_n705), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n816), .B(KEYINPUT99), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n493), .A2(new_n496), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT67), .B1(new_n492), .B2(new_n498), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n857));
  OAI211_X1 g432(.A(KEYINPUT98), .B(new_n505), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT98), .B1(new_n503), .B2(new_n505), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n853), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n850), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n629), .B(new_n480), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G162), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n850), .A2(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT103), .B(G37), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n868), .B(new_n869), .C1(new_n873), .C2(new_n866), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(new_n607), .B(G299), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n836), .B(new_n614), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n876), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n881), .ZN(new_n884));
  XOR2_X1   g459(.A(G305), .B(G288), .Z(new_n885));
  XNOR2_X1  g460(.A(G303), .B(G290), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G868), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(G868), .B2(new_n828), .ZN(G295));
  OAI21_X1  g466(.A(new_n890), .B1(G868), .B2(new_n828), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  XNOR2_X1  g469(.A(G168), .B(G301), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n836), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT106), .B1(new_n836), .B2(new_n895), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n876), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n836), .A2(new_n895), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(KEYINPUT105), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n836), .A2(new_n902), .A3(new_n895), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n880), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(KEYINPUT107), .A3(new_n887), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n887), .A2(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n899), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n876), .A2(new_n879), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(KEYINPUT108), .C1(new_n877), .C2(new_n876), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT108), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n898), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n883), .B1(new_n901), .B2(new_n903), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n887), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n887), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n899), .A2(new_n919), .A3(new_n904), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n918), .A2(KEYINPUT43), .A3(new_n869), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n894), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n918), .A2(new_n911), .A3(new_n869), .A4(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n894), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n893), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n922), .A2(new_n929), .A3(KEYINPUT109), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(G397));
  OAI21_X1  g506(.A(new_n505), .B1(new_n856), .B2(new_n857), .ZN(new_n932));
  AOI21_X1  g507(.A(G1384), .B1(new_n932), .B2(new_n855), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT50), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT112), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n936), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(G160), .A2(G40), .ZN(new_n939));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n861), .A2(new_n934), .A3(new_n940), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n742), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n861), .B2(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(G160), .A2(G40), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT117), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n933), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT117), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT98), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n858), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n952), .B2(new_n855), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n949), .B(new_n939), .C1(new_n953), .C2(KEYINPUT45), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n945), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1966), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n942), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G168), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n959), .A2(KEYINPUT51), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(new_n942), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT121), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT121), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n965), .B(new_n942), .C1(new_n955), .C2(new_n956), .ZN(new_n966));
  OAI21_X1  g541(.A(G8), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT122), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT122), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(G8), .C1(new_n964), .C2(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(new_n960), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n961), .B1(new_n972), .B2(KEYINPUT51), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n960), .B1(new_n964), .B2(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT62), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT62), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n960), .B1(new_n967), .B2(KEYINPUT122), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(new_n970), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n977), .B(new_n974), .C1(new_n980), .C2(new_n961), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n946), .A2(new_n947), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n939), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n751), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n944), .B1(new_n934), .B2(new_n933), .ZN(new_n986));
  INV_X1    g561(.A(G2090), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n986), .B(new_n987), .C1(new_n953), .C2(new_n934), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n958), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G166), .A2(new_n958), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n993));
  OAI22_X1  g568(.A1(G166), .A2(new_n958), .B1(KEYINPUT113), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n938), .A2(new_n941), .A3(new_n987), .A4(new_n939), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n958), .B(new_n995), .C1(new_n985), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G288), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(KEYINPUT52), .C1(G288), .C2(new_n1001), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n861), .A2(new_n939), .A3(new_n940), .ZN(new_n1008));
  OR2_X1    g583(.A1(G288), .A2(new_n1001), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(G8), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n547), .A2(G86), .ZN(new_n1011));
  INV_X1    g586(.A(new_n588), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1011), .B(new_n594), .C1(new_n1012), .C2(new_n586), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n589), .A2(new_n590), .A3(new_n1015), .A4(new_n594), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1014), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT49), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1008), .A3(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n958), .B1(new_n953), .B2(new_n939), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1003), .B1(new_n1022), .B2(new_n1009), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n997), .A2(new_n1000), .A3(KEYINPUT125), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT125), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n989), .B2(new_n996), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n999), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n938), .A2(new_n941), .A3(new_n939), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n938), .A2(new_n941), .A3(new_n1032), .A4(new_n939), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n716), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n984), .B2(G2078), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(G2078), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(new_n1036), .C1(new_n955), .C2(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1029), .A2(G171), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n976), .A2(new_n981), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1024), .B(KEYINPUT115), .Z(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n999), .ZN(new_n1043));
  AOI211_X1 g618(.A(G1976), .B(G288), .C1(new_n1022), .C2(new_n1019), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1016), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1022), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1043), .A2(KEYINPUT116), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n957), .A2(new_n958), .A3(G286), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n958), .B1(new_n985), .B2(new_n998), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(new_n996), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1000), .A2(KEYINPUT63), .ZN(new_n1052));
  AND4_X1   g627(.A1(new_n1042), .A2(new_n1049), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1054));
  NOR2_X1   g629(.A1(new_n1027), .A2(new_n999), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1049), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1047), .A2(new_n1048), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n955), .A2(new_n1038), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(G301), .A3(new_n1036), .A4(new_n1034), .ZN(new_n1059));
  INV_X1    g634(.A(new_n947), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n953), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(new_n939), .A3(new_n1037), .A4(new_n982), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1036), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1034), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1031), .A2(KEYINPUT123), .A3(new_n716), .A4(new_n1033), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT54), .B(new_n1059), .C1(new_n1067), .C2(G301), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1063), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(G301), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1039), .A2(G171), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT54), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1029), .B(new_n1068), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n934), .B1(new_n861), .B2(new_n940), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n939), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n798), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G299), .B(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n982), .A2(new_n939), .A3(new_n983), .A4(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1348), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1031), .A2(new_n1084), .A3(new_n1033), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n953), .A2(new_n818), .A3(new_n939), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n607), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1080), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1080), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(KEYINPUT61), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n982), .A2(new_n1098), .A3(new_n939), .A4(new_n983), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1008), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n550), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1095), .A2(new_n1097), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1085), .A2(KEYINPUT60), .A3(new_n1086), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1085), .A2(new_n1108), .A3(KEYINPUT60), .A4(new_n1086), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1087), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n607), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1105), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1107), .A2(new_n1112), .A3(new_n607), .A4(new_n1109), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1092), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1075), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n974), .B1(new_n980), .B2(new_n961), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1057), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1041), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n816), .B(new_n818), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n851), .B2(G1996), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n692), .B2(G1996), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n782), .A2(new_n786), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n781), .A2(new_n785), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G290), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n771), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT111), .Z(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(G1986), .B2(G290), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1061), .A2(new_n944), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1098), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT46), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1134), .B1(new_n851), .B2(new_n1123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT47), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1128), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1134), .A2(new_n1131), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1142), .A2(new_n1134), .B1(KEYINPUT48), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(KEYINPUT48), .B2(new_n1144), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1127), .B(KEYINPUT126), .Z(new_n1147));
  OAI22_X1  g722(.A1(new_n1125), .A2(new_n1147), .B1(G2067), .B2(new_n816), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1134), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1136), .A2(KEYINPUT127), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1135), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1041), .B2(new_n1120), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1155), .B2(new_n1150), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g732(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n874), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


