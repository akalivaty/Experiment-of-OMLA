//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G137), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT65), .B(G131), .Z(new_n197));
  AOI21_X1  g011(.A(new_n189), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G131), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n199), .A2(KEYINPUT66), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  OAI22_X1  g016(.A1(new_n198), .A2(new_n201), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT0), .B(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT66), .B1(new_n199), .B2(new_n200), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT11), .B1(new_n193), .B2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n193), .A2(G134), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n197), .A3(new_n189), .A4(new_n194), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n193), .A2(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n195), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n215), .A2(new_n219), .B1(G131), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(new_n210), .A3(KEYINPUT70), .A4(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n205), .ZN(new_n232));
  OAI21_X1  g046(.A(G128), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n210), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n214), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT71), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n241), .A2(new_n243), .A3(G116), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT72), .B1(new_n240), .B2(G116), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n239), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(new_n243), .A3(G116), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n248), .A4(new_n245), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n250), .A2(KEYINPUT73), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT73), .B1(new_n250), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT28), .B1(new_n238), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n214), .A3(new_n259), .A4(new_n237), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n212), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n209), .B(KEYINPUT64), .C1(new_n210), .C2(new_n211), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n203), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n215), .A2(new_n219), .B1(G131), .B2(new_n199), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n264), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n221), .A2(G131), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n198), .B2(new_n201), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n236), .B1(new_n222), .B2(new_n273), .ZN(new_n274));
  OAI22_X1  g088(.A1(new_n266), .A2(new_n269), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n258), .A2(new_n260), .B1(new_n275), .B2(new_n257), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT27), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n237), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n222), .A2(new_n273), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n226), .A2(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n271), .B2(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n203), .A2(new_n265), .A3(new_n261), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT67), .B1(new_n267), .B2(new_n268), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n284), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n257), .B(new_n283), .C1(new_n289), .C2(KEYINPUT30), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n281), .B1(new_n238), .B2(new_n257), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n290), .A2(new_n296), .A3(new_n291), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n282), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n237), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT30), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n275), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n301), .B2(new_n257), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT74), .B1(new_n302), .B2(new_n291), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n293), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT31), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n188), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n310), .B(new_n188), .C1(new_n298), .C2(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n238), .A2(new_n257), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n301), .B2(new_n257), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n315), .B2(new_n281), .ZN(new_n316));
  INV_X1    g130(.A(new_n314), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n290), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n281), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n276), .B2(new_n281), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n258), .A2(new_n260), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n238), .A2(new_n257), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n281), .A2(KEYINPUT29), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT77), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n329), .A3(new_n324), .A4(new_n325), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n312), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n309), .A2(new_n311), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G217), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(G234), .B2(new_n328), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT71), .B(G119), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G128), .ZN(new_n342));
  INV_X1    g156(.A(G128), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n240), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(new_n340), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G110), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT24), .B(G110), .Z(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT16), .ZN(new_n350));
  INV_X1    g164(.A(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(G125), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n204), .ZN(new_n358));
  OAI211_X1 g172(.A(G146), .B(new_n352), .C1(new_n356), .C2(new_n350), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT78), .B1(new_n356), .B2(G146), .ZN(new_n363));
  XNOR2_X1  g177(.A(G125), .B(G140), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n204), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n359), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n345), .A2(new_n348), .ZN(new_n369));
  INV_X1    g183(.A(G110), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n342), .C1(new_n345), .C2(new_n340), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n339), .B1(new_n362), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n359), .A3(new_n367), .ZN(new_n375));
  INV_X1    g189(.A(new_n339), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n361), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n328), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n335), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n383), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n373), .A2(new_n377), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n335), .A2(G902), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT80), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT81), .Z(new_n390));
  AND3_X1   g204(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n333), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  XNOR2_X1  g208(.A(G104), .B(G107), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT83), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(G101), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G104), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(G107), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n398), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(G104), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n404), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(G101), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n397), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n403), .A2(new_n401), .A3(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(new_n405), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT4), .B1(new_n413), .B2(G101), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n213), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n204), .A2(G143), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT1), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n210), .B2(G128), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n226), .B2(new_n230), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n397), .A2(new_n405), .A3(new_n409), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n411), .A2(new_n417), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n425), .A2(new_n203), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n411), .A2(new_n424), .A3(new_n417), .A4(new_n267), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n337), .A2(G227), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n429), .B(new_n430), .Z(new_n431));
  NOR3_X1   g245(.A1(new_n426), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n236), .A2(new_n410), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n422), .A2(new_n423), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n203), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT12), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT84), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  INV_X1    g252(.A(new_n421), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n231), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n410), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n285), .A2(new_n423), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n267), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n443), .B2(KEYINPUT12), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(KEYINPUT12), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n427), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n432), .B1(new_n447), .B2(new_n431), .ZN(new_n448));
  OAI21_X1  g262(.A(G469), .B1(new_n448), .B2(G902), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n431), .B1(new_n426), .B2(new_n428), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n428), .A2(new_n431), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n431), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n425), .A2(new_n203), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(new_n427), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT85), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G469), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n328), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G221), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT9), .B(G234), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(new_n328), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n394), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT86), .B(new_n466), .C1(new_n449), .C2(new_n461), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  INV_X1    g285(.A(G122), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT98), .B(KEYINPUT14), .C1(new_n472), .C2(G116), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(G116), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n247), .A2(G122), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n474), .C1(KEYINPUT14), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT98), .B1(new_n475), .B2(KEYINPUT14), .ZN(new_n477));
  OAI21_X1  g291(.A(G107), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT97), .ZN(new_n479));
  XNOR2_X1  g293(.A(G116), .B(G122), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n400), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n479), .A2(new_n474), .A3(new_n475), .A4(new_n400), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n206), .A2(G128), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n343), .A2(G143), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT96), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT96), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n487), .A2(new_n488), .A3(new_n191), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G134), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n478), .B(new_n483), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n191), .B1(new_n487), .B2(new_n488), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n480), .B(new_n400), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT13), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(G134), .C1(KEYINPUT13), .C2(new_n484), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n464), .A2(new_n334), .A3(G953), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n494), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n328), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n471), .B1(new_n503), .B2(KEYINPUT99), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT99), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(new_n328), .C1(new_n501), .C2(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(new_n508), .B2(new_n471), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n277), .A2(G143), .A3(G214), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G143), .B1(new_n277), .B2(G214), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT18), .B(G131), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n337), .A3(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n206), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n364), .A2(new_n204), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n363), .B2(new_n366), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n365), .B1(new_n364), .B2(new_n204), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n365), .A2(new_n353), .A3(new_n355), .A4(new_n204), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n524), .A2(new_n525), .B1(new_n204), .B2(new_n364), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n519), .A4(new_n514), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n402), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n197), .A2(new_n517), .A3(new_n511), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n197), .A2(new_n517), .A3(KEYINPUT94), .A4(new_n511), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n200), .B1(new_n512), .B2(new_n513), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n358), .A2(new_n359), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n537), .A2(new_n535), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n529), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n531), .B1(new_n529), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n328), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G475), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n356), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n364), .A2(KEYINPUT19), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n204), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT19), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT19), .B1(new_n353), .B2(new_n355), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT95), .B(new_n204), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n554), .A2(new_n555), .A3(new_n359), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n531), .B1(new_n529), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n546), .B(new_n547), .C1(new_n542), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n529), .A2(new_n531), .A3(new_n541), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n359), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT95), .B1(new_n551), .B2(new_n204), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n555), .A2(new_n566), .B1(new_n523), .B2(new_n528), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n563), .B1(new_n567), .B2(new_n531), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n546), .B1(new_n568), .B2(new_n547), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n545), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n337), .A2(G952), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(G234), .B2(G237), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n328), .B(new_n337), .C1(G234), .C2(G237), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT21), .B(G898), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n510), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G214), .B1(G237), .B2(G902), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n254), .A2(new_n255), .B1(new_n415), .B2(new_n416), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT89), .ZN(new_n580));
  INV_X1    g394(.A(G113), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n244), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n252), .A2(new_n248), .A3(new_n245), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n582), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n580), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n583), .B(KEYINPUT89), .C1(new_n585), .C2(new_n582), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n253), .A3(new_n410), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n590));
  OAI221_X1 g404(.A(new_n590), .B1(new_n415), .B2(new_n416), .C1(new_n254), .C2(new_n255), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n579), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(G110), .B(G122), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n579), .A2(new_n595), .A3(new_n591), .A4(new_n589), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(KEYINPUT6), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT6), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n598), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n213), .A2(G125), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n285), .B2(G125), .ZN(new_n601));
  INV_X1    g415(.A(G224), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT7), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(KEYINPUT91), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n607), .B2(new_n603), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n593), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT5), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n585), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n253), .B1(new_n584), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(new_n410), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n587), .A2(new_n253), .A3(new_n588), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n410), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n601), .A2(KEYINPUT91), .A3(KEYINPUT7), .A4(new_n604), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n609), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n619), .B2(new_n596), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(G210), .B1(G237), .B2(G902), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(KEYINPUT92), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n623), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n606), .B2(new_n620), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n576), .B(new_n577), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n468), .A2(new_n469), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n393), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(new_n398), .Z(G3));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n631));
  INV_X1    g445(.A(new_n432), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n436), .B(new_n267), .C1(new_n441), .C2(new_n442), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n435), .A2(new_n436), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n438), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n428), .B1(new_n635), .B2(new_n437), .ZN(new_n636));
  OAI211_X1 g450(.A(G469), .B(new_n632), .C1(new_n636), .C2(new_n455), .ZN(new_n637));
  NAND2_X1  g451(.A1(G469), .A2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n446), .A2(new_n453), .B1(new_n457), .B2(KEYINPUT85), .ZN(new_n640));
  AOI211_X1 g454(.A(G469), .B(G902), .C1(new_n640), .C2(new_n452), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n467), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n462), .A2(new_n394), .A3(new_n467), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n391), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n282), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n296), .B1(new_n302), .B2(new_n291), .ZN(new_n647));
  INV_X1    g461(.A(new_n297), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n305), .B1(new_n304), .B2(KEYINPUT31), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT74), .B(new_n291), .C1(new_n290), .C2(new_n293), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n187), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n298), .B2(new_n307), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(new_n312), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n631), .B1(new_n645), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n655), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n468), .A2(new_n469), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT100), .A4(new_n391), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n621), .A2(new_n622), .ZN(new_n661));
  INV_X1    g475(.A(new_n622), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n606), .A2(new_n662), .A3(new_n620), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n661), .A2(new_n577), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n570), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n503), .A2(new_n470), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT101), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n503), .A2(new_n668), .A3(new_n470), .ZN(new_n669));
  OR3_X1    g483(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT33), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT33), .B1(new_n501), .B2(new_n502), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n470), .A2(G902), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n667), .A2(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n665), .A2(new_n674), .A3(new_n575), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n660), .A2(new_n664), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NOR3_X1   g492(.A1(new_n570), .A2(new_n509), .A3(new_n575), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n660), .A2(new_n664), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NOR2_X1   g496(.A1(new_n655), .A2(new_n627), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n375), .A2(new_n361), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n388), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n384), .A2(new_n385), .A3(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n468), .A2(new_n469), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n573), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n572), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n570), .A2(new_n509), .A3(new_n697), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n577), .A2(new_n661), .A3(new_n663), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n384), .A2(new_n385), .A3(new_n687), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n643), .A2(new_n699), .A3(new_n644), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n333), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n343), .ZN(G30));
  XNOR2_X1  g517(.A(new_n696), .B(KEYINPUT39), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n658), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT40), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n653), .A2(new_n310), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n315), .A2(new_n319), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n317), .A2(new_n319), .A3(new_n324), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n328), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n624), .A2(new_n626), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT38), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n665), .A2(new_n509), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n577), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n715), .A2(new_n700), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n706), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  INV_X1    g534(.A(new_n332), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n707), .A2(new_n708), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n665), .A2(new_n674), .A3(new_n697), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n661), .A2(new_n577), .A3(new_n663), .ZN(new_n726));
  INV_X1    g540(.A(new_n723), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n689), .A2(new_n722), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI21_X1  g544(.A(new_n460), .B1(new_n459), .B2(new_n328), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n467), .A3(new_n461), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n726), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n722), .A2(new_n391), .A3(new_n675), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  AND2_X1   g551(.A1(new_n722), .A2(new_n734), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n391), .A2(new_n679), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT103), .B(G116), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G18));
  AND2_X1   g556(.A1(new_n700), .A2(new_n576), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  AOI21_X1  g559(.A(new_n281), .B1(new_n323), .B2(new_n324), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(KEYINPUT31), .B2(new_n304), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n647), .B2(new_n648), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n187), .B(KEYINPUT104), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n391), .B(new_n750), .C1(new_n312), .C2(new_n654), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n716), .A2(new_n661), .A3(new_n577), .A4(new_n663), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n733), .A3(new_n575), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  NOR2_X1   g570(.A1(new_n641), .A2(new_n731), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n664), .A2(new_n467), .A3(new_n723), .A4(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n700), .B(new_n750), .C1(new_n654), .C2(new_n312), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n354), .ZN(G27));
  NAND2_X1  g575(.A1(new_n322), .A2(new_n331), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n308), .A2(KEYINPUT32), .B1(new_n762), .B2(G472), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n653), .A2(new_n764), .A3(new_n310), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT105), .B1(new_n308), .B2(KEYINPUT32), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n577), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n624), .A2(new_n768), .A3(new_n626), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n466), .B1(new_n449), .B2(new_n461), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n769), .A2(new_n770), .A3(new_n723), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n391), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT42), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n769), .A2(new_n770), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n722), .A2(new_n774), .A3(new_n775), .A4(new_n391), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n202), .ZN(G33));
  NAND4_X1  g592(.A1(new_n722), .A2(new_n774), .A3(new_n391), .A4(new_n698), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n665), .B1(new_n674), .B2(KEYINPUT106), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n674), .A2(KEYINPUT106), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n570), .A2(new_n674), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n785), .A2(KEYINPUT107), .B1(KEYINPUT43), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n655), .A3(new_n700), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT44), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n448), .A2(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n448), .A2(KEYINPUT45), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n638), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n641), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n467), .A3(new_n704), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(new_n769), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT108), .B(G137), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G39));
  AND3_X1   g617(.A1(new_n799), .A2(KEYINPUT47), .A3(new_n467), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT47), .B1(new_n799), .B2(new_n467), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n333), .A2(new_n392), .A3(new_n723), .A4(new_n769), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  OR2_X1    g623(.A1(G952), .A2(G953), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n695), .B1(new_n786), .B2(new_n789), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n752), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n734), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n571), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n769), .A2(new_n467), .A3(new_n757), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n811), .A2(new_n391), .A3(new_n767), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n392), .A2(new_n695), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n665), .A2(new_n674), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n816), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n665), .A3(new_n674), .A4(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(new_n759), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n811), .A2(new_n829), .A3(new_n817), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n467), .A2(new_n715), .A3(new_n768), .A4(new_n757), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n812), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT50), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n757), .A2(new_n466), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n806), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n812), .A2(new_n769), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n827), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n838), .B1(new_n806), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT113), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n843), .B1(new_n848), .B2(new_n837), .ZN(new_n849));
  AOI211_X1 g663(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n836), .C2(new_n847), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT117), .B(new_n842), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n333), .A2(new_n701), .B1(new_n759), .B2(new_n758), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT109), .ZN(new_n857));
  INV_X1    g671(.A(new_n753), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n642), .A2(new_n700), .A3(new_n697), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n713), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n733), .A2(new_n727), .A3(new_n726), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n829), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n862), .B(new_n863), .C1(new_n333), .C2(new_n701), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n857), .A2(new_n729), .A3(new_n860), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  INV_X1    g680(.A(new_n701), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n760), .B1(new_n867), .B2(new_n722), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n729), .A4(new_n860), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT110), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n866), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n722), .A2(new_n391), .A3(new_n774), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n875), .A2(new_n775), .B1(new_n772), .B2(KEYINPUT42), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n722), .B(new_n734), .C1(new_n739), .C2(new_n743), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n735), .A3(new_n755), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n510), .A2(new_n570), .A3(new_n697), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n769), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n689), .A2(new_n722), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n771), .A2(new_n829), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(new_n779), .A3(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n393), .A2(new_n628), .B1(new_n689), .B2(new_n683), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n824), .B1(new_n665), .B2(new_n510), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n888), .A2(new_n714), .A3(new_n575), .A4(new_n768), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n656), .A2(new_n659), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT53), .A4(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n880), .A2(new_n881), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n872), .A2(new_n874), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n876), .A2(new_n879), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n886), .A2(new_n887), .A3(new_n890), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n658), .A2(new_n700), .A3(new_n724), .A4(new_n728), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n860), .B1(new_n898), .B2(new_n333), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT52), .B1(new_n899), .B2(new_n856), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT111), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(new_n870), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n900), .B2(new_n870), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n897), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n894), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n872), .A2(new_n874), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(new_n905), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n911), .B2(new_n894), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n810), .B1(new_n855), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n757), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(KEYINPUT49), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n391), .A2(new_n467), .A3(new_n577), .A4(new_n788), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(KEYINPUT49), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n820), .A3(new_n715), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(new_n919), .ZN(G75));
  NAND2_X1  g734(.A1(new_n597), .A2(new_n599), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT118), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT55), .Z(new_n923));
  INV_X1    g737(.A(new_n605), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n328), .B1(new_n893), .B2(new_n906), .ZN(new_n925));
  AOI211_X1 g739(.A(KEYINPUT56), .B(new_n924), .C1(new_n925), .C2(G210), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n893), .A2(new_n906), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(G210), .A3(G902), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n605), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n337), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n926), .A2(new_n930), .A3(new_n923), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G51));
  NAND2_X1  g750(.A1(new_n907), .A2(KEYINPUT119), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n893), .A2(new_n906), .A3(new_n938), .A4(new_n894), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n927), .A2(KEYINPUT54), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n638), .B(KEYINPUT57), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n459), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n925), .A2(G469), .A3(new_n794), .A4(new_n793), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n568), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n932), .ZN(G60));
  XNOR2_X1  g765(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n470), .A2(new_n328), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n912), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n672), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n954), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n932), .B1(new_n941), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI211_X1 g776(.A(KEYINPUT121), .B(new_n932), .C1(new_n941), .C2(new_n959), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G63));
  XNOR2_X1  g778(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n334), .A2(new_n328), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n927), .A2(new_n686), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n927), .A2(new_n967), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n933), .B(new_n968), .C1(new_n969), .C2(new_n386), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n574), .B2(new_n602), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n879), .A2(new_n890), .A3(new_n887), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n922), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(G898), .B2(new_n337), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  AOI21_X1  g792(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n301), .B(new_n551), .Z(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(G900), .B2(G953), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n800), .A2(new_n391), .A3(new_n858), .A4(new_n767), .ZN(new_n982));
  AND4_X1   g796(.A1(new_n779), .A2(new_n808), .A3(new_n801), .A4(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n857), .A2(new_n729), .A3(new_n864), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n876), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n981), .B1(new_n985), .B2(G953), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n979), .B1(new_n986), .B2(KEYINPUT125), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n888), .B(KEYINPUT124), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n393), .A2(new_n988), .A3(new_n705), .A4(new_n769), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n808), .A2(new_n801), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n719), .A2(new_n984), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n719), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n980), .B1(new_n995), .B2(G953), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n986), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n987), .B(new_n997), .Z(G72));
  NAND3_X1  g812(.A1(new_n316), .A2(new_n304), .A3(new_n320), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1001), .ZN(new_n1003));
  INV_X1    g817(.A(new_n985), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n974), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n315), .A2(new_n319), .ZN(new_n1006));
  OAI221_X1 g820(.A(new_n933), .B1(new_n911), .B2(new_n1002), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n995), .B2(new_n974), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n709), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1009), .A2(new_n1013), .A3(new_n709), .A4(new_n1010), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1012), .B2(new_n1014), .ZN(G57));
endmodule


