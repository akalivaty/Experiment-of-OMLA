//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G97), .A2(G257), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n202), .B1(new_n247), .B2(G20), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n252), .A2(new_n253), .B1(new_n202), .B2(new_n249), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G150), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n211), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(G20), .B2(new_n203), .ZN(new_n260));
  INV_X1    g0060(.A(new_n251), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(KEYINPUT9), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(KEYINPUT9), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n266), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n266), .A2(KEYINPUT68), .A3(G222), .A4(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  AND2_X1   g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n284), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(G200), .B1(new_n280), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n280), .A2(new_n289), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n265), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n280), .A2(new_n289), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G190), .B1(new_n263), .B2(new_n264), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(KEYINPUT71), .A3(KEYINPUT10), .A4(new_n290), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n279), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n273), .B2(new_n287), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n308), .A2(new_n309), .A3(new_n272), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n301), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n286), .ZN(new_n312));
  INV_X1    g0112(.A(new_n288), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(G238), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G200), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n269), .B2(new_n258), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n251), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT11), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n248), .A2(G68), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT12), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n327), .C2(new_n326), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n247), .A2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n252), .A2(G68), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n316), .A2(G190), .A3(new_n318), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n320), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n319), .A2(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n316), .A2(G179), .A3(new_n318), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(new_n318), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n317), .B1(new_n311), .B2(new_n314), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(G169), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n338), .B1(new_n346), .B2(new_n334), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n297), .A2(KEYINPUT69), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n291), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n291), .A2(G179), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n349), .B(new_n262), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G238), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n267), .A2(new_n355), .B1(new_n356), .B2(new_n266), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n308), .A2(new_n309), .A3(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n301), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n312), .B1(G244), .B2(new_n313), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n361), .A2(G169), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(KEYINPUT70), .ZN(new_n364));
  INV_X1    g0164(.A(G87), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(KEYINPUT15), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(KEYINPUT15), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n257), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n261), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n252), .A2(G77), .A3(new_n332), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G77), .B2(new_n248), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n361), .A2(new_n348), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n362), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n359), .A2(G190), .A3(new_n360), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n361), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n300), .A2(new_n347), .A3(new_n354), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n390));
  INV_X1    g0190(.A(new_n252), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n373), .A2(new_n332), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n248), .B2(new_n373), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n266), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G68), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n321), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n255), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n261), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n397), .B2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT16), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n393), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n266), .A2(G226), .A3(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT73), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n411), .B(new_n413), .C1(new_n273), .C2(new_n268), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n301), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n286), .B1(new_n309), .B2(new_n288), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT74), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n286), .B(new_n419), .C1(new_n309), .C2(new_n288), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n414), .B2(new_n301), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n416), .A2(new_n421), .B1(new_n422), .B2(G200), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n390), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n321), .B1(new_n395), .B2(new_n396), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n406), .B1(new_n425), .B2(new_n403), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n409), .A2(new_n251), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n393), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AND4_X1   g0230(.A1(new_n427), .A2(new_n423), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT76), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n428), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  INV_X1    g0234(.A(new_n421), .ZN(new_n435));
  AOI21_X1  g0235(.A(G179), .B1(new_n414), .B2(new_n301), .ZN(new_n436));
  INV_X1    g0236(.A(new_n417), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n415), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n435), .A2(new_n436), .B1(new_n438), .B2(new_n351), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n433), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n433), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n423), .A2(new_n427), .A3(new_n428), .ZN(new_n443));
  INV_X1    g0243(.A(new_n390), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n410), .A2(new_n423), .A3(new_n430), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n432), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n389), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n305), .A2(new_n307), .A3(G257), .A4(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(new_n272), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G294), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(new_n301), .ZN(new_n455));
  INV_X1    g0255(.A(G41), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n247), .B(G45), .C1(new_n456), .C2(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n247), .A4(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n459), .A2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n462), .A3(new_n283), .A4(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(new_n279), .C1(new_n457), .C2(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n455), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n454), .A2(new_n301), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n466), .A4(new_n465), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(G169), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n455), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G179), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n247), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n252), .A2(G107), .A3(new_n477), .ZN(new_n478));
  OR3_X1    g0278(.A1(new_n248), .A2(KEYINPUT25), .A3(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT25), .B1(new_n248), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(KEYINPUT80), .A3(new_n479), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n356), .A3(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT78), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n211), .A2(G107), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT79), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT78), .B(KEYINPUT23), .C1(new_n211), .C2(G107), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n489), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n488), .A3(new_n487), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n356), .A2(G20), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT78), .B1(new_n497), .B2(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT79), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n266), .A2(new_n211), .A3(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n266), .A2(new_n502), .A3(new_n211), .A4(G87), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n495), .A2(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n251), .B1(new_n504), .B2(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n503), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n506), .A2(KEYINPUT24), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n485), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n472), .A2(new_n510), .A3(new_n474), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n476), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n507), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n504), .A2(KEYINPUT24), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n251), .ZN(new_n517));
  AOI21_X1  g0317(.A(G190), .B1(new_n468), .B2(new_n471), .ZN(new_n518));
  INV_X1    g0318(.A(new_n467), .ZN(new_n519));
  AOI21_X1  g0319(.A(G200), .B1(new_n519), .B2(new_n469), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n517), .B(new_n485), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(G1698), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n305), .A2(new_n307), .A3(G238), .A4(new_n272), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n301), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  INV_X1    g0328(.A(G45), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G1), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n247), .A2(new_n281), .A3(G45), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n279), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n211), .B1(new_n302), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n365), .A2(new_n538), .A3(new_n356), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n305), .A2(new_n307), .A3(new_n211), .A4(G68), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n258), .B2(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n251), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n249), .B1(new_n364), .B2(new_n369), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n252), .A2(G87), .A3(new_n477), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n532), .B1(new_n526), .B2(new_n301), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n535), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n364), .A2(new_n369), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n252), .A2(new_n477), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n544), .B(new_n545), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n548), .A2(new_n351), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n348), .B(new_n532), .C1(new_n526), .C2(new_n301), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(G1698), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(new_n272), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n301), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n279), .C1(new_n457), .C2(new_n463), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n465), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n351), .ZN(new_n567));
  INV_X1    g0367(.A(new_n565), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n561), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n558), .A4(new_n559), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n571), .B2(new_n301), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n348), .A3(new_n465), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n255), .A2(G77), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n575), .A2(new_n538), .A3(G107), .ZN(new_n576));
  XNOR2_X1  g0376(.A(G97), .B(G107), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n575), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n574), .B1(new_n578), .B2(new_n211), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n356), .B1(new_n395), .B2(new_n396), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n251), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n248), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n552), .B2(new_n538), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n567), .A2(new_n573), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n581), .A2(new_n585), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n566), .A2(G200), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n572), .A2(G190), .A3(new_n465), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n557), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n252), .A2(G116), .A3(new_n477), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n249), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n250), .A2(new_n210), .B1(G20), .B2(new_n594), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n558), .B(new_n211), .C1(G33), .C2(new_n538), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n593), .B(new_n595), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n305), .A2(new_n307), .A3(G264), .A4(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n305), .A2(new_n307), .A3(G257), .A4(new_n272), .ZN(new_n602));
  INV_X1    g0402(.A(G303), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n266), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n301), .ZN(new_n605));
  OAI211_X1 g0405(.A(G270), .B(new_n279), .C1(new_n457), .C2(new_n463), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n465), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n600), .B1(new_n607), .B2(G200), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n292), .B2(new_n607), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(G169), .A3(new_n600), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n465), .A2(new_n606), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n600), .A2(G179), .A3(new_n605), .A4(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n607), .A2(KEYINPUT21), .A3(G169), .A4(new_n600), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n609), .A2(new_n612), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n592), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n450), .A2(new_n522), .A3(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n354), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n346), .A2(new_n334), .B1(new_n337), .B2(new_n382), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n432), .A2(new_n448), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n442), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(new_n300), .ZN(new_n623));
  INV_X1    g0423(.A(new_n450), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n468), .A2(new_n471), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n520), .B1(new_n625), .B2(new_n292), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n509), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n591), .A2(new_n587), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n517), .A2(new_n485), .B1(new_n472), .B2(new_n474), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT84), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n553), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT83), .B1(new_n554), .B2(new_n555), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n527), .A2(G179), .A3(new_n533), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(new_n351), .C2(new_n548), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n550), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n475), .A2(new_n509), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n615), .A2(new_n614), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n351), .B1(new_n613), .B2(new_n605), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT21), .B1(new_n643), .B2(new_n600), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT84), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n629), .A2(new_n632), .A3(new_n640), .A4(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n566), .A2(new_n351), .B1(new_n581), .B2(new_n585), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n573), .A3(new_n556), .A4(new_n550), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n638), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n634), .A2(new_n637), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n553), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n567), .A2(new_n573), .A3(new_n586), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n550), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n623), .B1(new_n624), .B2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n247), .A2(new_n211), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n509), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n512), .A2(new_n521), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n666), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n512), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n600), .A2(new_n666), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n631), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n616), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n645), .A2(new_n666), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n522), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n630), .A2(new_n669), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n676), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n207), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n539), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n214), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n617), .A2(new_n521), .A3(new_n512), .A4(new_n669), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n519), .A2(new_n469), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n534), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n613), .A2(G179), .A3(new_n605), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT85), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT30), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n691), .A2(new_n693), .A3(new_n572), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n473), .A2(new_n572), .A3(new_n548), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n695), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n548), .A2(G179), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n607), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n700), .B2(new_n607), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n566), .A2(new_n690), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n697), .B(new_n699), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n666), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT87), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT87), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n712), .B(KEYINPUT31), .C1(new_n706), .C2(new_n666), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n591), .A2(new_n587), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n640), .A3(new_n521), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n512), .B2(new_n645), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n654), .A2(new_n557), .A3(new_n655), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n638), .A2(new_n587), .A3(new_n639), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n653), .B(new_n720), .C1(new_n721), .C2(new_n655), .ZN(new_n722));
  OAI211_X1 g0522(.A(KEYINPUT29), .B(new_n669), .C1(new_n719), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n666), .B1(new_n648), .B2(new_n657), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n716), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n688), .B1(new_n726), .B2(G1), .ZN(G364));
  AND2_X1   g0527(.A1(new_n211), .A2(G13), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n247), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n683), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n210), .B1(G20), .B2(new_n351), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n211), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n292), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n356), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n308), .B(new_n737), .C1(G87), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT90), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT89), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT32), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT32), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n292), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n211), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n538), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n742), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n752), .A2(new_n385), .A3(G190), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n755), .A2(G77), .B1(G68), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n753), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n385), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n757), .B1(new_n202), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n758), .A2(G200), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n751), .B(new_n761), .C1(G58), .C2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n741), .A2(new_n747), .A3(new_n748), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n762), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n766), .B1(new_n736), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n750), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(G294), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n756), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n772), .B1(new_n754), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n743), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n266), .B(new_n774), .C1(G329), .C2(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G326), .A2(new_n759), .B1(new_n739), .B2(G303), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n734), .B1(new_n764), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n733), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n682), .A2(new_n308), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n594), .B2(new_n682), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n245), .A2(G45), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT88), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n682), .A2(new_n266), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n215), .B2(G45), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n732), .B(new_n779), .C1(new_n783), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n782), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n674), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n731), .B1(new_n674), .B2(G330), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G330), .B2(new_n674), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  OAI22_X1  g0597(.A1(new_n384), .A2(new_n386), .B1(new_n378), .B2(new_n669), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n381), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n362), .A2(new_n379), .A3(new_n380), .A4(new_n669), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n724), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n731), .B1(new_n803), .B2(new_n716), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n716), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n733), .A2(new_n780), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n731), .B1(G77), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT91), .Z(new_n809));
  OAI21_X1  g0609(.A(new_n308), .B1(new_n738), .B2(new_n356), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT92), .Z(new_n811));
  OAI22_X1  g0611(.A1(new_n743), .A2(new_n773), .B1(new_n754), .B2(new_n594), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G283), .B2(new_n756), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n751), .B1(G303), .B2(new_n759), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n736), .A2(new_n365), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G294), .B2(new_n762), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n755), .A2(G159), .B1(G150), .B2(new_n756), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n765), .B2(new_n819), .C1(new_n820), .C2(new_n760), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n266), .B1(new_n743), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G50), .B2(new_n739), .ZN(new_n826));
  INV_X1    g0626(.A(new_n736), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n769), .A2(G58), .B1(new_n827), .B2(G68), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n821), .A2(new_n822), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n817), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n809), .B1(new_n831), .B2(new_n733), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n802), .B2(new_n781), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n805), .A2(new_n833), .ZN(G384));
  NAND2_X1  g0634(.A1(new_n577), .A2(new_n575), .ZN(new_n835));
  INV_X1    g0635(.A(new_n576), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n838), .A2(new_n839), .A3(new_n594), .A4(new_n213), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT36), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n400), .A2(new_n214), .A3(new_n269), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n202), .A2(G68), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n247), .B(G13), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT96), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n334), .B(new_n666), .C1(new_n346), .C2(new_n338), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n345), .A2(new_n341), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n342), .B1(new_n319), .B2(G169), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n334), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n334), .A2(new_n666), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n337), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n666), .B(new_n801), .C1(new_n648), .C2(new_n657), .ZN(new_n854));
  INV_X1    g0654(.A(new_n800), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n664), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n251), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT93), .B1(new_n426), .B2(new_n251), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n425), .A2(new_n406), .A3(new_n403), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n861), .B2(new_n393), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n449), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT94), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n251), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT93), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n251), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n393), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n443), .B1(new_n870), .B2(new_n664), .ZN(new_n871));
  INV_X1    g0671(.A(new_n439), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n865), .B(KEYINPUT37), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n433), .A2(new_n439), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n664), .B(KEYINPUT95), .Z(new_n876));
  NAND2_X1  g0676(.A1(new_n433), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n877), .A3(new_n443), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n439), .B1(new_n861), .B2(new_n393), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n862), .A2(new_n881), .A3(new_n443), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n865), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT38), .B(new_n864), .C1(new_n880), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n864), .B1(new_n880), .B2(new_n883), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n856), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n442), .A2(new_n876), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n846), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n853), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n658), .A2(new_n669), .A3(new_n802), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n800), .ZN(new_n893));
  INV_X1    g0693(.A(new_n884), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n871), .B2(new_n873), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT94), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n879), .A3(new_n874), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n897), .B2(new_n864), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n893), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n889), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT96), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n878), .B(KEYINPUT37), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n445), .A2(new_n446), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n877), .B1(new_n442), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n886), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n884), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n346), .A2(new_n334), .A3(new_n669), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n902), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n890), .A2(new_n901), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n623), .B1(new_n624), .B2(new_n725), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n801), .B1(new_n847), .B2(new_n852), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n709), .A2(new_n710), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n689), .A2(new_n917), .A3(new_n707), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n916), .A2(KEYINPUT40), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n887), .B2(new_n884), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n922), .B2(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n450), .A2(new_n918), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(G330), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n247), .B2(new_n728), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n915), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n845), .B1(new_n929), .B2(new_n930), .ZN(G367));
  INV_X1    g0731(.A(new_n788), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n783), .B1(new_n238), .B2(new_n932), .C1(new_n207), .C2(new_n551), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n731), .ZN(new_n934));
  INV_X1    g0734(.A(G150), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n819), .A2(new_n760), .B1(new_n765), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G58), .B2(new_n739), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n771), .A2(new_n744), .B1(new_n754), .B2(new_n202), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n308), .B(new_n938), .C1(G137), .C2(new_n775), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n736), .A2(new_n269), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G68), .B2(new_n769), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n769), .A2(G107), .B1(new_n759), .B2(G311), .ZN(new_n943));
  AOI22_X1  g0743(.A1(G303), .A2(new_n762), .B1(new_n827), .B2(G97), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n266), .B1(G294), .B2(new_n756), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G317), .A2(new_n775), .B1(new_n755), .B2(G283), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT100), .B1(new_n739), .B2(G116), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT46), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n942), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n547), .A2(new_n669), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n653), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n640), .B2(new_n952), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT97), .Z(new_n955));
  OAI221_X1 g0755(.A(new_n934), .B1(new_n734), .B2(new_n951), .C1(new_n955), .C2(new_n792), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n717), .B1(new_n588), .B2(new_n669), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n587), .B2(new_n669), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n680), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT45), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT44), .B1(new_n680), .B2(new_n959), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n680), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(new_n676), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n678), .B1(new_n670), .B2(new_n677), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(new_n675), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n726), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n965), .B(new_n969), .C1(KEYINPUT99), .C2(new_n676), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n964), .A2(new_n676), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT99), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n726), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n683), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n730), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n959), .A2(new_n678), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT42), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n587), .B1(new_n957), .B2(new_n512), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n669), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT98), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT98), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n979), .A2(new_n982), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n955), .B(KEYINPUT43), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n671), .A2(new_n675), .A3(new_n959), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n988), .B(new_n989), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n956), .B1(new_n977), .B2(new_n990), .ZN(G387));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n969), .B2(new_n684), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n968), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n726), .C2(new_n967), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n257), .A2(G50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT103), .B(KEYINPUT50), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n685), .ZN(new_n999));
  AOI211_X1 g0799(.A(G45), .B(new_n999), .C1(G68), .C2(G77), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1001), .B2(KEYINPUT102), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT102), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n788), .B1(new_n529), .B2(new_n235), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n784), .A2(new_n999), .B1(new_n356), .B2(new_n682), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT101), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n732), .B1(new_n1008), .B2(new_n783), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n308), .B1(new_n775), .B2(G150), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n269), .B2(new_n738), .C1(new_n538), .C2(new_n736), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT104), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n771), .A2(new_n257), .B1(new_n754), .B2(new_n321), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT105), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n370), .A2(new_n769), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n762), .B1(new_n759), .B2(G159), .ZN(new_n1016));
  AND4_X1   g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n769), .A2(G283), .B1(new_n739), .B2(G294), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n755), .A2(G303), .B1(G311), .B2(new_n756), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n762), .A2(G317), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n766), .C2(new_n760), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT106), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT49), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n266), .B1(new_n775), .B2(G326), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n594), .B2(new_n736), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1025), .B2(KEYINPUT49), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1017), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1009), .B1(new_n1030), .B2(new_n734), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n671), .B2(new_n782), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n967), .B2(new_n730), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n995), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT108), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n995), .A2(KEYINPUT108), .A3(new_n1033), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(G393));
  AND2_X1   g0838(.A1(new_n965), .A2(new_n971), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n730), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G150), .A2(new_n759), .B1(new_n762), .B2(G159), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT51), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n771), .A2(new_n202), .B1(new_n754), .B2(new_n257), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n308), .B(new_n1043), .C1(G143), .C2(new_n775), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n750), .A2(new_n269), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n815), .B(new_n1045), .C1(G68), .C2(new_n739), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n762), .B1(new_n759), .B2(G317), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT52), .Z(new_n1049));
  INV_X1    g0849(.A(G294), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n743), .A2(new_n766), .B1(new_n754), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n266), .B(new_n1051), .C1(G303), .C2(new_n756), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n738), .A2(new_n767), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n737), .B(new_n1053), .C1(G116), .C2(new_n769), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n734), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n783), .B1(new_n538), .B2(new_n207), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n242), .B2(new_n788), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n732), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n958), .B2(new_n792), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1040), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1039), .A2(new_n969), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n684), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n970), .A2(new_n973), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(G390));
  NAND2_X1  g0866(.A1(new_n902), .A2(new_n909), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n892), .A2(new_n800), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n911), .B1(new_n1068), .B2(new_n853), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G330), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n708), .B2(new_n714), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n802), .A3(new_n853), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n669), .B(new_n799), .C1(new_n719), .C2(new_n722), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n800), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n853), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n910), .A3(new_n907), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1071), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n918), .A2(G330), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1080), .A2(new_n916), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1069), .B1(new_n902), .B2(new_n909), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1078), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n450), .A2(new_n1080), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n623), .C1(new_n624), .C2(new_n725), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n853), .B1(new_n1073), .B2(new_n802), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1068), .B1(new_n1087), .B2(new_n1081), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n918), .A2(G330), .A3(new_n802), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1076), .B1(new_n891), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1074), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1086), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1079), .A2(new_n1084), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n683), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT109), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1092), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1093), .A2(KEYINPUT109), .A3(new_n683), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1079), .A2(new_n1084), .A3(new_n730), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1067), .A2(new_n780), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n731), .B1(new_n373), .B2(new_n807), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT110), .Z(new_n1105));
  OAI22_X1  g0905(.A1(new_n594), .A2(new_n765), .B1(new_n760), .B2(new_n767), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1045), .B(new_n1106), .C1(G68), .C2(new_n827), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n308), .B1(new_n743), .B2(new_n1050), .C1(new_n365), .C2(new_n738), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT111), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n771), .A2(new_n356), .B1(new_n754), .B2(new_n538), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1107), .B(new_n1111), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n771), .A2(new_n820), .B1(new_n754), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n308), .B(new_n1114), .C1(G125), .C2(new_n775), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n738), .A2(new_n935), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G132), .A2(new_n762), .B1(new_n827), .B2(G50), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n769), .A2(G159), .B1(new_n759), .B2(G128), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1103), .B(new_n1105), .C1(new_n734), .C2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1102), .A2(KEYINPUT112), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT112), .B1(new_n1102), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT113), .B1(new_n1101), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1101), .A2(new_n1125), .A3(KEYINPUT113), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(G378));
  AOI21_X1  g0929(.A(KEYINPUT96), .B1(new_n899), .B2(new_n900), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n902), .A2(new_n909), .A3(new_n911), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n354), .A2(new_n296), .A3(new_n299), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n262), .A2(new_n857), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT55), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n354), .A2(new_n296), .A3(new_n1140), .A4(new_n299), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1136), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1134), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1138), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1136), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1133), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1072), .B1(new_n907), .B2(new_n919), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n922), .C2(KEYINPUT40), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n887), .A2(new_n884), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n921), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT40), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n920), .A2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1132), .A2(new_n901), .A3(new_n1151), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1151), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n913), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1158), .A2(new_n1160), .A3(KEYINPUT118), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT118), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n730), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n769), .A2(G150), .B1(new_n759), .B2(G125), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n765), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n738), .A2(new_n1113), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n771), .A2(new_n824), .B1(new_n754), .B2(new_n820), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT59), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(G33), .A2(G41), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT114), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n736), .A2(new_n744), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G124), .C2(new_n775), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n765), .A2(new_n356), .B1(new_n736), .B2(new_n399), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n759), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n456), .B(new_n308), .C1(new_n743), .C2(new_n767), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n750), .A2(new_n321), .B1(new_n738), .B2(new_n269), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G97), .C2(new_n756), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n551), .C2(new_n754), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1174), .B(new_n202), .C1(G41), .C2(new_n266), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1177), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n733), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT115), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n732), .B(new_n1190), .C1(new_n202), .C2(new_n806), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1149), .B2(new_n781), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1163), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1086), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1093), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT119), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n683), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1196), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT118), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1132), .A2(new_n901), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1159), .A2(new_n913), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1158), .A2(new_n1160), .A3(KEYINPUT118), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1200), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1206), .B2(KEYINPUT57), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n684), .B1(new_n1209), .B2(new_n1196), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n1198), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1193), .B1(new_n1207), .B2(new_n1211), .ZN(G375));
  AND2_X1   g1012(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1086), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n976), .A3(new_n1098), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n853), .A2(new_n781), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT120), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n732), .B1(new_n321), .B2(new_n806), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n771), .A2(new_n594), .B1(new_n743), .B2(new_n603), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n266), .B(new_n1219), .C1(G107), .C2(new_n755), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n940), .B1(G97), .B2(new_n739), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G283), .A2(new_n762), .B1(new_n759), .B2(G294), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n1015), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n769), .A2(G50), .B1(new_n762), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n744), .B2(new_n738), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n266), .B1(new_n771), .B2(new_n1113), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n743), .A2(new_n1165), .B1(new_n754), .B2(new_n935), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n760), .A2(new_n824), .B1(new_n736), .B2(new_n399), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT122), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n734), .B1(new_n1232), .B2(KEYINPUT122), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1217), .B(new_n1218), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1213), .B2(new_n729), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1215), .A2(new_n1238), .ZN(G381));
  NAND2_X1  g1039(.A1(new_n1163), .A2(new_n1192), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1196), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1241), .A2(new_n1208), .B1(new_n1210), .B2(new_n1198), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1211), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT123), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1065), .B(new_n956), .C1(new_n977), .C2(new_n990), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1036), .A2(new_n796), .A3(new_n1037), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G384), .A2(new_n1246), .A3(G381), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1102), .A2(new_n1122), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1101), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OR3_X1    g1052(.A1(new_n1245), .A2(new_n1248), .A3(new_n1252), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n665), .A2(G213), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT124), .Z(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(new_n1245), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(new_n1194), .A2(new_n730), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1192), .B(new_n1258), .C1(new_n1241), .C2(new_n975), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1251), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1101), .A2(KEYINPUT113), .A3(new_n1125), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1126), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(G375), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1255), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1098), .A2(KEYINPUT60), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1265), .A2(new_n1214), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n683), .B1(new_n1265), .B2(new_n1214), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1238), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1238), .B(new_n1269), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1263), .A2(new_n1264), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1255), .A2(G2897), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1275), .B(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1244), .A2(G378), .B1(new_n1251), .B2(new_n1259), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1255), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1263), .A2(new_n1284), .A3(new_n1264), .A4(new_n1276), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1278), .A2(new_n1279), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n796), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1289), .B2(new_n1247), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1247), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1291), .A2(new_n1288), .A3(KEYINPUT126), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G390), .A2(G387), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1246), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1288), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1287), .A3(new_n1247), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1293), .A2(new_n1296), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1295), .A2(new_n1299), .A3(new_n1298), .A4(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1286), .A2(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1264), .A4(new_n1276), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1281), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1277), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1251), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1262), .B2(G375), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(new_n1275), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1305), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1314), .B(new_n1276), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1303), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(G402));
endmodule


