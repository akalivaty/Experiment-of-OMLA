//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(KEYINPUT3), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n462), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(new_n470), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n469), .A2(new_n462), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n462), .A2(new_n464), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n485), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n487), .A2(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n462), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n490), .A2(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT67), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT67), .A2(G651), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT6), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT68), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n498), .A2(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT69), .B(G88), .Z(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n498), .B2(new_n500), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n496), .A2(new_n497), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n503), .B2(new_n505), .ZN(new_n514));
  AND2_X1   g089(.A1(G75), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(new_n510), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n506), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n503), .A2(new_n505), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n521), .A2(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(G168));
  NAND2_X1  g102(.A1(new_n521), .A2(G64), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n512), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n509), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n506), .A2(G90), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  NAND2_X1  g110(.A1(new_n506), .A2(G81), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n509), .A2(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n536), .B(new_n537), .C1(new_n511), .C2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n521), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(G65), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G91), .B2(new_n506), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n509), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT67), .A2(G651), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(G49), .B(G543), .C1(new_n565), .C2(new_n499), .ZN(new_n566));
  OAI211_X1 g141(.A(G87), .B(new_n521), .C1(new_n565), .C2(new_n499), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT74), .A4(new_n568), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n503), .B2(new_n505), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n512), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(G86), .B(new_n521), .C1(new_n565), .C2(new_n499), .ZN(new_n578));
  OAI211_X1 g153(.A(G48), .B(G543), .C1(new_n565), .C2(new_n499), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(G85), .A2(new_n506), .B1(new_n509), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n511), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n506), .A2(G92), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n586), .B(KEYINPUT76), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n552), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n472), .A2(new_n488), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(G2100), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n477), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n479), .A2(G123), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT78), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT17), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2084), .B(G2090), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n640), .B2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  INV_X1    g221(.A(new_n642), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n647), .A2(new_n643), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n644), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n655), .A2(new_n660), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n660), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n659), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G23), .B(new_n569), .S(G16), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT80), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT33), .B(G1976), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G22), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G166), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n677), .A2(new_n678), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n477), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n479), .A2(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n470), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(G1986), .Z(new_n699));
  NAND4_X1  g274(.A1(new_n688), .A2(new_n689), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT81), .B(KEYINPUT36), .Z(new_n701));
  NOR3_X1   g276(.A1(new_n700), .A2(KEYINPUT82), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n477), .A2(G139), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT25), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n705), .C1(new_n470), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G33), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G2072), .Z(new_n709));
  INV_X1    g284(.A(KEYINPUT24), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(G34), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n474), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2084), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G28), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n618), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n718), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT84), .Z(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT29), .B(G2090), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n718), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n477), .A2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n479), .A2(G128), .ZN(new_n732));
  OR2_X1    g307(.A1(G104), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(new_n718), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2067), .ZN(new_n738));
  NOR4_X1   g313(.A1(new_n716), .A2(new_n724), .A3(new_n728), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n679), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n543), .B2(new_n679), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1341), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n679), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n479), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI22_X1  g329(.A1(G105), .A2(new_n472), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n749), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G32), .B(new_n756), .S(G29), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n679), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n679), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1961), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n758), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2078), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n759), .A2(new_n762), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n679), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n679), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1966), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n761), .A2(G1961), .B1(G2078), .B2(new_n765), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G4), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n597), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT83), .B(G1348), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n739), .A2(new_n748), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n702), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n700), .A2(KEYINPUT36), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(KEYINPUT82), .C1(new_n700), .C2(new_n701), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(G311));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(G150));
  XOR2_X1   g359(.A(KEYINPUT88), .B(G860), .Z(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n604), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT38), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT86), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n790), .A2(new_n791), .A3(new_n511), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n790), .B2(new_n511), .ZN(new_n793));
  AOI22_X1  g368(.A1(G93), .A2(new_n506), .B1(new_n509), .B2(G55), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT87), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n792), .A2(new_n794), .A3(KEYINPUT87), .A4(new_n793), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n797), .A2(new_n539), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n541), .A2(new_n542), .A3(new_n795), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n789), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n786), .B1(new_n803), .B2(KEYINPUT39), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(KEYINPUT39), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n797), .A2(new_n798), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n786), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT37), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(G145));
  NAND2_X1  g384(.A1(new_n477), .A2(G142), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n479), .A2(G130), .ZN(new_n812));
  OR2_X1    g387(.A1(G106), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n694), .B(KEYINPUT92), .ZN(new_n818));
  INV_X1    g393(.A(new_n611), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n694), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n611), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n611), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n818), .A2(new_n819), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(new_n826), .A3(new_n816), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n824), .A2(KEYINPUT93), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n707), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n756), .ZN(new_n835));
  INV_X1    g410(.A(G164), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n735), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n736), .A3(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n832), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n830), .A2(new_n842), .A3(new_n840), .A4(new_n831), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT94), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n474), .B(KEYINPUT89), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n722), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n830), .A2(new_n831), .B1(new_n842), .B2(new_n840), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(G37), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n849), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n840), .A2(new_n842), .A3(new_n828), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT95), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n840), .A2(new_n842), .A3(new_n858), .A4(new_n828), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n855), .A2(new_n860), .A3(KEYINPUT96), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT96), .B1(new_n855), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g439(.A(new_n606), .B(new_n801), .Z(new_n865));
  AND2_X1   g440(.A1(new_n787), .A2(G299), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n787), .A2(G299), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n866), .B2(new_n867), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n787), .A2(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n787), .A2(G299), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n870), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  XOR2_X1   g454(.A(G290), .B(new_n569), .Z(new_n880));
  XOR2_X1   g455(.A(G303), .B(G305), .Z(new_n881));
  XOR2_X1   g456(.A(new_n880), .B(new_n881), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n806), .A2(new_n600), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  INV_X1    g465(.A(new_n882), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n892));
  NAND3_X1  g467(.A1(G171), .A2(G168), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G168), .B1(KEYINPUT97), .B2(G301), .ZN(new_n894));
  NAND2_X1  g469(.A1(G171), .A2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n801), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n893), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n800), .A3(new_n799), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n868), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n800), .B2(new_n799), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n898), .A2(KEYINPUT98), .A3(new_n800), .A4(new_n799), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n891), .B(new_n900), .C1(new_n905), .C2(new_n876), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT100), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(KEYINPUT100), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n900), .B1(new_n905), .B2(new_n876), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n911), .B2(new_n882), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g489(.A(KEYINPUT99), .B(G37), .C1(new_n911), .C2(new_n882), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n909), .B(new_n910), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n903), .A2(new_n904), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n868), .A3(new_n897), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n897), .A2(new_n899), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n876), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n920), .B2(new_n882), .ZN(new_n921));
  INV_X1    g496(.A(new_n908), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n906), .A2(KEYINPUT100), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n890), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT43), .B1(new_n907), .B2(new_n908), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n927), .A2(KEYINPUT43), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n890), .B2(new_n929), .ZN(G397));
  INV_X1    g505(.A(G2067), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n735), .B(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n756), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n696), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n694), .A2(new_n936), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n935), .A2(new_n937), .B1(G2067), .B2(new_n735), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n490), .B2(new_n494), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n466), .A2(G40), .A3(new_n471), .A4(new_n473), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n932), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n946), .B2(new_n756), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n933), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  NOR2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n694), .A2(new_n936), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n932), .A2(new_n934), .A3(new_n937), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n944), .B2(new_n959), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n945), .B(new_n952), .C1(new_n956), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n943), .B1(new_n940), .B2(KEYINPUT50), .ZN(new_n962));
  INV_X1    g537(.A(G2090), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(new_n939), .C1(new_n490), .C2(new_n494), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n943), .B1(new_n940), .B2(new_n941), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT45), .B(new_n939), .C1(new_n490), .C2(new_n494), .ZN(new_n968));
  AOI21_X1  g543(.A(G1971), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT55), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(G303), .A2(G8), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(KEYINPUT55), .ZN(new_n977));
  AOI22_X1  g552(.A1(G303), .A2(G8), .B1(new_n977), .B2(new_n974), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(G303), .A2(G8), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n977), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT102), .A3(new_n975), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n970), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g561(.A1(G305), .A2(G1981), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  NAND3_X1  g567(.A1(G305), .A2(KEYINPUT104), .A3(G1981), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n940), .B2(new_n943), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n488), .A2(new_n489), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n491), .A2(new_n493), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n943), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n566), .A2(new_n567), .A3(G1976), .A4(new_n568), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT103), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n571), .A2(new_n1010), .A3(new_n572), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1005), .A2(new_n1008), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1006), .B(KEYINPUT103), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT52), .B1(new_n1013), .B2(new_n996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n986), .B1(new_n997), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n991), .A2(new_n993), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT49), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1005), .A3(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(KEYINPUT109), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n985), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(G2084), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n962), .A2(new_n965), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1966), .B1(new_n967), .B2(new_n968), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1027), .A2(new_n998), .A3(G286), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT107), .B(new_n1004), .C1(new_n1003), .C2(new_n964), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n965), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT108), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n1033));
  INV_X1    g608(.A(new_n965), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n962), .B2(KEYINPUT107), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1037), .A3(new_n963), .ZN(new_n1038));
  INV_X1    g613(.A(new_n969), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n998), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n976), .A2(new_n978), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1022), .B(new_n1028), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1028), .A2(KEYINPUT63), .ZN(new_n1046));
  INV_X1    g621(.A(new_n985), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT105), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n997), .B2(new_n1015), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1020), .A2(KEYINPUT105), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n970), .A2(new_n1041), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1046), .A2(new_n1047), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G288), .A2(G1976), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n994), .B2(new_n995), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n996), .B1(new_n1056), .B2(new_n990), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT106), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1051), .A2(new_n985), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT106), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1057), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1045), .A2(new_n1053), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1027), .A2(G168), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n942), .A2(new_n1004), .A3(new_n968), .ZN(new_n1065));
  OAI211_X1 g640(.A(G168), .B(new_n1024), .C1(new_n1065), .C2(G1966), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT51), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1022), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1022), .B(KEYINPUT122), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n942), .A2(new_n1076), .A3(new_n1004), .A4(new_n968), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT119), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n967), .A2(new_n1079), .A3(new_n1076), .A4(new_n968), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n962), .A2(new_n965), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1077), .A2(new_n1088), .A3(new_n1082), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1081), .A2(new_n1084), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1070), .B2(KEYINPUT62), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .A4(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n555), .B2(new_n557), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n555), .A2(new_n557), .A3(new_n1094), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1956), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n967), .A2(new_n968), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n746), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n555), .A2(new_n557), .A3(new_n1094), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1095), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1101), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1098), .B(KEYINPUT118), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1348), .B1(new_n962), .B2(new_n965), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n940), .A2(G2067), .A3(new_n943), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n597), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n940), .B2(new_n943), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT115), .B(G1996), .Z(new_n1122));
  NAND4_X1  g697(.A1(new_n942), .A2(new_n1004), .A3(new_n968), .A4(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT116), .B(new_n1118), .C1(new_n940), .C2(new_n943), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1125), .A2(new_n543), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1125), .B2(new_n543), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1117), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1115), .A2(new_n787), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n597), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1116), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT113), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1103), .A2(new_n1136), .A3(new_n1106), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1096), .A2(new_n1138), .A3(new_n1097), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT114), .B1(new_n1104), .B2(new_n1095), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1101), .B1(new_n1143), .B2(new_n746), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1110), .B1(new_n1144), .B2(new_n1105), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1112), .A2(new_n1134), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1132), .B(KEYINPUT112), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1107), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT121), .B(G2078), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1065), .A2(KEYINPUT53), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1091), .B1(G171), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1155), .A2(new_n1156), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(KEYINPUT124), .A3(new_n1153), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n1161));
  AOI21_X1  g736(.A(G301), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1156), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1159), .A2(KEYINPUT123), .A3(G301), .A4(new_n1081), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1090), .B2(G171), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1074), .A2(new_n1168), .A3(new_n1075), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1063), .B(new_n1093), .C1(new_n1158), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  XNOR2_X1  g746(.A(G290), .B(G1986), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n944), .B1(new_n959), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n961), .B1(new_n1174), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(G319), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G227), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n637), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1180), .A2(KEYINPUT126), .ZN(new_n1181));
  OR2_X1    g755(.A1(new_n1180), .A2(KEYINPUT126), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n671), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n863), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n929), .ZN(G308));
  OR2_X1    g759(.A1(new_n1184), .A2(new_n929), .ZN(G225));
endmodule


