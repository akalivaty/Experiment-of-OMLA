//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n463), .A2(new_n461), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  OR2_X1    g049(.A1(new_n474), .A2(new_n465), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n469), .A2(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n470), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n473), .A2(G138), .A3(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n486), .A2(KEYINPUT69), .A3(new_n488), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g078(.A(new_n503), .B(KEYINPUT70), .Z(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n506), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n504), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(new_n502), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n505), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n522), .A2(G51), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n520), .B2(new_n521), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n500), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  NAND3_X1  g109(.A1(new_n506), .A2(new_n508), .A3(G64), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(new_n521), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(new_n500), .A3(G90), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G52), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n522), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(KEYINPUT72), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n511), .A2(new_n546), .B1(new_n513), .B2(new_n541), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n502), .B1(new_n535), .B2(new_n536), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n544), .A2(new_n549), .ZN(G171));
  NAND3_X1  g125(.A1(new_n506), .A2(new_n508), .A3(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(KEYINPUT73), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n555), .A2(G651), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n511), .A2(new_n558), .B1(new_n513), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n506), .A2(new_n508), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n511), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n572), .A2(G651), .B1(new_n573), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n522), .A2(G53), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n522), .A2(KEYINPUT9), .A3(G53), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(G299));
  AND2_X1   g154(.A1(new_n544), .A2(new_n549), .ZN(G301));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  OAI21_X1  g156(.A(G89), .B1(new_n509), .B2(new_n510), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n570), .B1(new_n582), .B2(new_n530), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n524), .A2(new_n526), .ZN(new_n584));
  OAI211_X1 g159(.A(G51), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G286));
  NAND2_X1  g164(.A1(new_n573), .A2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n522), .A2(G49), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n522), .A2(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n511), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n502), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n502), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT75), .Z(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n511), .A2(new_n604), .B1(new_n513), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OR3_X1    g184(.A1(new_n511), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n570), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n522), .A2(G54), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT10), .B1(new_n511), .B2(new_n609), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n610), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G171), .B2(new_n618), .ZN(G284));
  XOR2_X1   g195(.A(G284), .B(KEYINPUT76), .Z(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(new_n617), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  OAI21_X1  g203(.A(KEYINPUT77), .B1(new_n562), .B2(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  MUX2_X1   g206(.A(KEYINPUT77), .B(new_n629), .S(new_n631), .Z(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g208(.A(new_n479), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n634), .A2(KEYINPUT78), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n470), .A2(G135), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT78), .B1(new_n634), .B2(new_n635), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n636), .A2(new_n637), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2100), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT80), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2451), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT81), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT82), .Z(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT83), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n670), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(new_n668), .A3(new_n665), .ZN(new_n674));
  INV_X1    g249(.A(new_n668), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n665), .A3(new_n666), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT85), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n691), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT87), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT86), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n696), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G5), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G171), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G1961), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT101), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n704), .A2(G20), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G299), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1956), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n641), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G26), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT96), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n479), .A2(G128), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n470), .A2(G140), .ZN(new_n720));
  NOR2_X1   g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2067), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G29), .A2(G32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n470), .A2(G141), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT100), .Z(new_n729));
  AND3_X1   g304(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT26), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n730), .B(new_n732), .C1(new_n479), .C2(G129), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT27), .B(G1996), .Z(new_n737));
  AOI211_X1 g312(.A(new_n715), .B(new_n726), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n714), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n714), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT29), .Z(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n714), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n714), .ZN(new_n745));
  INV_X1    g320(.A(G2078), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n748), .A2(new_n714), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G160), .B2(new_n714), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n738), .A2(new_n743), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n741), .A2(new_n742), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n562), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G16), .B2(G19), .ZN(new_n757));
  INV_X1    g332(.A(G1341), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n704), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n704), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(G28), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n765), .A2(new_n766), .A3(new_n714), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n755), .A2(new_n759), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n706), .B2(G1961), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n736), .A2(new_n737), .B1(new_n758), .B2(new_n757), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n754), .A2(new_n768), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n773));
  MUX2_X1   g348(.A(G6), .B(G305), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT32), .B(G1981), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n704), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n704), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n777), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G24), .ZN(new_n795));
  XOR2_X1   g370(.A(G290), .B(KEYINPUT91), .Z(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT92), .B(G1986), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n714), .A2(G25), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n479), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n470), .A2(G131), .ZN(new_n803));
  OR2_X1    g378(.A1(G95), .A2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n804), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT89), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n800), .B(new_n801), .C1(new_n807), .C2(G29), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n800), .B2(new_n801), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT90), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n799), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n773), .B1(new_n794), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g390(.A(KEYINPUT36), .B(new_n813), .C1(new_n792), .C2(new_n793), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n708), .B(new_n772), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n626), .A2(G16), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G4), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT95), .B(G1348), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(G29), .A2(G33), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  INV_X1    g398(.A(G139), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n466), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n470), .A2(KEYINPUT97), .A3(G139), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT25), .Z(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n473), .A2(G127), .ZN(new_n833));
  NAND2_X1  g408(.A1(G115), .A2(G2104), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n465), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n822), .B1(new_n837), .B2(new_n714), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT99), .B(G2072), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n817), .A2(new_n821), .A3(new_n840), .ZN(G311));
  INV_X1    g416(.A(new_n772), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n794), .A2(new_n814), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n794), .A2(new_n773), .A3(new_n814), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n821), .ZN(new_n847));
  INV_X1    g422(.A(new_n840), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n708), .ZN(G150));
  NAND3_X1  g424(.A1(new_n506), .A2(new_n508), .A3(G67), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G651), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n522), .A2(G55), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n539), .A2(new_n500), .A3(G93), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n511), .A2(new_n858), .B1(new_n513), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n502), .B1(new_n850), .B2(new_n851), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT103), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT105), .B(G860), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n626), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n862), .A2(new_n857), .B1(new_n557), .B2(new_n561), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n855), .B(new_n856), .C1(new_n871), .C2(new_n502), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n557), .A2(new_n561), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT104), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(G145));
  NAND4_X1  g455(.A1(new_n492), .A2(new_n486), .A3(new_n495), .A4(new_n488), .ZN(new_n881));
  NAND2_X1  g456(.A1(G160), .A2(new_n484), .ZN(new_n882));
  INV_X1    g457(.A(new_n641), .ZN(new_n883));
  INV_X1    g458(.A(new_n476), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n468), .B2(new_n471), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n484), .B1(new_n885), .B2(new_n475), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n477), .A2(G162), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n641), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n881), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n881), .A3(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n807), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n837), .A2(new_n644), .ZN(new_n895));
  INV_X1    g470(.A(new_n644), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n832), .A2(new_n896), .A3(new_n836), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n832), .B2(new_n836), .ZN(new_n899));
  AOI211_X1 g474(.A(new_n644), .B(new_n835), .C1(new_n830), .C2(new_n831), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n900), .A3(new_n807), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n892), .B(new_n893), .C1(new_n898), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n894), .A3(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n807), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(new_n893), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n891), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n479), .A2(G130), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n470), .A2(G142), .ZN(new_n909));
  NOR2_X1   g484(.A1(G106), .A2(G2105), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n734), .B(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(new_n723), .Z(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n902), .A2(new_n906), .A3(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT106), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n916), .A2(new_n921), .A3(new_n917), .A4(new_n918), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(G395));
  XOR2_X1   g500(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n617), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G299), .A2(new_n617), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n874), .B(new_n630), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n937), .B(KEYINPUT108), .Z(new_n938));
  NOR2_X1   g513(.A1(new_n928), .A2(new_n929), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G305), .B(G288), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(G303), .ZN(new_n943));
  INV_X1    g518(.A(G290), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT109), .Z(new_n948));
  NOR2_X1   g523(.A1(new_n941), .A2(new_n946), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n618), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n948), .A2(new_n950), .B1(new_n618), .B2(new_n863), .ZN(G295));
  AOI22_X1  g526(.A1(new_n948), .A2(new_n950), .B1(new_n618), .B2(new_n863), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n544), .A2(new_n549), .A3(new_n533), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G301), .B2(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n874), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n587), .A2(new_n588), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G171), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n954), .C1(new_n873), .C2(new_n870), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n874), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n934), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n960), .A2(new_n934), .A3(KEYINPUT111), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n956), .A2(new_n939), .A3(new_n959), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT112), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n945), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n943), .B(G290), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n917), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n960), .A2(new_n962), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n956), .A2(new_n959), .B1(new_n939), .B2(new_n926), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n939), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(KEYINPUT41), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n945), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n973), .A2(new_n981), .A3(new_n982), .A4(new_n917), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n974), .A2(KEYINPUT43), .B1(new_n983), .B2(KEYINPUT113), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n953), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n973), .A2(new_n981), .A3(new_n917), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT114), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n973), .A2(new_n981), .A3(new_n988), .A4(new_n917), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n974), .A2(new_n982), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT44), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n985), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n985), .B2(new_n992), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(G397));
  XNOR2_X1  g571(.A(new_n723), .B(G2067), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n734), .B2(G1996), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n881), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(KEYINPUT45), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n472), .A2(G40), .A3(new_n475), .A4(new_n476), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1005), .B2(G1996), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1003), .A2(new_n1001), .A3(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(KEYINPUT116), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(new_n735), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n807), .A2(new_n810), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n807), .A2(new_n810), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1009), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G290), .B(G1986), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n498), .B2(new_n999), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(new_n885), .A3(G40), .A4(new_n475), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n780), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n498), .B2(new_n999), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n881), .A2(new_n1026), .A3(new_n999), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(new_n885), .A3(G40), .A4(new_n475), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(new_n1029), .A3(G2090), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1020), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n742), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n1024), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT55), .Z(new_n1036));
  NAND4_X1  g611(.A1(new_n1031), .A2(new_n1034), .A3(G8), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  OAI221_X1 g613(.A(G8), .B1(new_n1038), .B2(G288), .C1(new_n1003), .C2(new_n1000), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n596), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n599), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1045), .A2(G1981), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(G305), .B2(G1981), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1045), .A2(new_n1049), .A3(G1981), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT49), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1050), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1053), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1003), .A2(new_n1000), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1042), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n498), .A2(new_n1026), .A3(new_n999), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1004), .B(new_n1061), .C1(new_n1026), .C2(new_n1001), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1024), .B1(new_n1062), .B2(G2090), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1036), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n746), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1002), .A2(new_n1069), .A3(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1004), .A3(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1032), .A2(G1961), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1037), .A2(new_n1060), .A3(new_n1066), .A4(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G301), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1004), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n762), .B1(new_n1078), .B2(new_n1002), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1032), .A2(new_n752), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(G168), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1056), .A2(KEYINPUT123), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(G8), .A3(new_n533), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT62), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1084), .A2(new_n1086), .A3(new_n1091), .A4(new_n1088), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1077), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1021), .A2(new_n1023), .A3(G1996), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT58), .B(G1341), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1055), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n562), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n562), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1348), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1055), .A2(new_n725), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1105), .A2(new_n617), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n617), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n626), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1101), .A2(new_n1103), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n623), .B(KEYINPUT121), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT57), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1067), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1062), .A2(KEYINPUT120), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT120), .B1(new_n1062), .B2(new_n1118), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1115), .B(new_n1117), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1102), .A2(new_n1101), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1121), .C1(new_n617), .C2(new_n1110), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1037), .A2(new_n1060), .A3(new_n1066), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G301), .B(KEYINPUT54), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1023), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1071), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1070), .A2(new_n1133), .A3(new_n1074), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1075), .A2(new_n1131), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1130), .A2(new_n1089), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1093), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1031), .A2(G8), .A3(new_n1034), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1065), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1056), .B(G286), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1037), .A3(new_n1060), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1037), .A2(new_n1060), .A3(new_n1066), .A4(new_n1141), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1138), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1037), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1060), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1058), .A2(new_n1038), .A3(new_n783), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(G1981), .B2(G305), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1057), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1145), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1019), .B1(new_n1137), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n723), .A2(G2067), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1154));
  OR3_X1    g729(.A1(new_n1154), .A2(KEYINPUT124), .A3(new_n1005), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1005), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT48), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1155), .B(new_n1156), .C1(new_n1017), .C2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1012), .B(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n997), .A2(new_n734), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1162), .A2(new_n1009), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT126), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(new_n1166), .A3(new_n1163), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT47), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT47), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1165), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1159), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1152), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(G227), .ZN(new_n1175));
  AND3_X1   g749(.A1(new_n919), .A2(new_n1175), .A3(new_n702), .ZN(new_n1176));
  OR2_X1    g750(.A1(new_n975), .A2(new_n984), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n1176), .A2(G319), .A3(new_n663), .A4(new_n1177), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


