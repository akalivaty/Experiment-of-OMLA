//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G127gat), .A2(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G113gat), .B2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT67), .B(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n207), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(new_n212), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n205), .B(new_n206), .C1(new_n215), .C2(new_n209), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT2), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n217), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n213), .A2(new_n216), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n224), .A2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT76), .B1(new_n217), .B2(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n224), .A2(new_n234), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n224), .B2(new_n234), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT75), .B1(new_n246), .B2(new_n217), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(new_n229), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n234), .A3(new_n243), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(KEYINPUT75), .A3(new_n217), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n236), .B(new_n242), .C1(new_n247), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT39), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n241), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n217), .A2(new_n235), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(KEYINPUT80), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(KEYINPUT80), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G57gat), .ZN(new_n267));
  INV_X1    g066(.A(G85gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n258), .A3(new_n256), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT40), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n259), .A2(new_n260), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n256), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n217), .A2(new_n235), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n247), .B2(new_n253), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n238), .B1(new_n237), .B2(new_n239), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n217), .A2(new_n235), .A3(KEYINPUT76), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n255), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT5), .B(new_n275), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n250), .A2(new_n217), .A3(new_n251), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n252), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n287), .A2(new_n236), .A3(new_n242), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n269), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT26), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT26), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n294), .A3(new_n299), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n302), .A2(new_n308), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  OAI211_X1 g112(.A(G183gat), .B(G190gat), .C1(new_n313), .C2(KEYINPUT24), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(KEYINPUT65), .A3(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n321), .A3(new_n303), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT25), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n319), .A2(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n315), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n317), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n327), .A3(new_n328), .A4(new_n303), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n312), .A2(new_n323), .A3(new_n332), .A4(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n339));
  INV_X1    g138(.A(G197gat), .ZN(new_n340));
  INV_X1    g139(.A(G204gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G211gat), .A2(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n344), .B(new_n347), .C1(new_n338), .C2(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n335), .A2(new_n355), .A3(new_n336), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  INV_X1    g159(.A(G64gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G92gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n362), .B(G92gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n293), .B1(new_n359), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n335), .A2(new_n336), .A3(new_n355), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n355), .B1(new_n335), .B2(new_n336), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT30), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n379), .A3(new_n366), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n264), .A2(KEYINPUT40), .A3(new_n269), .A4(new_n270), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n273), .A2(new_n292), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n383), .A2(new_n292), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n271), .A2(new_n272), .B1(new_n376), .B2(new_n381), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT81), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n251), .A2(new_n333), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n355), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  INV_X1    g192(.A(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n348), .A2(new_n338), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n333), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n348), .A2(new_n338), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n243), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n235), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n392), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n349), .B2(new_n350), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n235), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n392), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(G22gat), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n405), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n395), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n402), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT31), .B(G50gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n403), .A2(new_n406), .A3(G22gat), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n410), .B1(new_n409), .B2(new_n402), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT79), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n413), .A3(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n371), .B2(new_n372), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n357), .A2(KEYINPUT37), .A3(new_n358), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n364), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n426), .A2(KEYINPUT38), .B1(new_n366), .B2(new_n359), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n290), .A2(KEYINPUT6), .A3(new_n291), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n283), .A2(new_n269), .A3(new_n289), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n269), .B1(new_n283), .B2(new_n289), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n427), .B(new_n428), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n369), .A2(KEYINPUT38), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n373), .B2(KEYINPUT37), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n425), .A2(KEYINPUT82), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n436), .B(KEYINPUT83), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n373), .A2(new_n437), .A3(KEYINPUT37), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n425), .A2(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT83), .B1(new_n444), .B2(new_n436), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n422), .B1(new_n434), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n390), .A2(new_n447), .A3(KEYINPUT84), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT84), .B1(new_n390), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n330), .A2(new_n237), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n312), .A2(new_n323), .A3(new_n217), .A4(new_n329), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  INV_X1    g253(.A(G227gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n394), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n456), .B(KEYINPUT64), .Z(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT70), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n460), .A3(new_n454), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n456), .B1(new_n451), .B2(new_n452), .ZN(new_n464));
  NOR2_X1   g263(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NOR4_X1   g269(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n468), .A4(new_n465), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n453), .A2(new_n457), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G71gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G99gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n462), .B(new_n474), .C1(new_n470), .C2(new_n471), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n476), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n476), .B2(new_n485), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n464), .ZN(new_n490));
  INV_X1    g289(.A(new_n465), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n469), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g292(.A(new_n471), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n474), .B1(new_n495), .B2(new_n462), .ZN(new_n496));
  INV_X1    g295(.A(new_n485), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n483), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n476), .A2(new_n484), .A3(new_n485), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT78), .ZN(new_n502));
  INV_X1    g301(.A(new_n428), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n290), .B2(new_n291), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT77), .B(new_n269), .C1(new_n283), .C2(new_n289), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND4_X1   g306(.A1(new_n287), .A2(new_n236), .A3(new_n242), .A4(new_n288), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT5), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n286), .A2(new_n252), .B1(KEYINPUT4), .B2(new_n276), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n256), .B1(new_n259), .B2(new_n202), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n508), .B1(new_n275), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT6), .B1(new_n513), .B2(new_n269), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n502), .B1(new_n515), .B2(new_n382), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT77), .B1(new_n513), .B2(new_n269), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n432), .A2(new_n504), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n428), .ZN(new_n520));
  INV_X1    g319(.A(new_n382), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n501), .B1(new_n523), .B2(new_n422), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n486), .A2(new_n422), .A3(new_n487), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n525), .A2(new_n521), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n450), .A2(new_n524), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G57gat), .B(G64gat), .Z(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  INV_X1    g332(.A(G78gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n480), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT86), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(KEYINPUT86), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n545), .A2(KEYINPUT86), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n541), .A2(new_n543), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n539), .A2(KEYINPUT21), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT91), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT19), .ZN(new_n552));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT20), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n554), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n536), .B(new_n537), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  AND3_X1   g362(.A1(new_n555), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n555), .B2(new_n556), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G162gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G29gat), .ZN(new_n570));
  INV_X1    g369(.A(G36gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT14), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(new_n570), .B2(new_n571), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT15), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n572), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n573), .B2(new_n572), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G43gat), .B(G50gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n576), .B2(KEYINPUT15), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n583), .B1(new_n577), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT17), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT93), .B1(new_n592), .B2(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n593), .A2(new_n596), .A3(KEYINPUT93), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n268), .B2(new_n363), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n591), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n590), .A2(new_n587), .ZN(new_n613));
  INV_X1    g412(.A(new_n609), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n607), .A2(new_n608), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(G134gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(G134gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n569), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n568), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n566), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n531), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n613), .A2(new_n546), .A3(new_n549), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n546), .A2(new_n549), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n590), .B2(new_n587), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n589), .A2(new_n591), .A3(new_n635), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT87), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n642), .A3(new_n634), .A4(new_n638), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT88), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT18), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n634), .A3(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n647), .B2(KEYINPUT88), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n640), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G197gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT11), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n304), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n640), .B(new_n655), .C1(new_n645), .C2(new_n649), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n557), .B1(new_n614), .B2(new_n615), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n539), .A2(new_n606), .A3(new_n609), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n539), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT94), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT95), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n305), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n341), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n663), .A2(new_n665), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n662), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n670), .A2(new_n671), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n666), .A2(new_n667), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n669), .B1(new_n679), .B2(new_n661), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT94), .B(new_n662), .C1(new_n666), .C2(new_n667), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n675), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT95), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n677), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n674), .B1(new_n685), .B2(new_n668), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n660), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n633), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n520), .B(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT97), .B(G1gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1324gat));
  OAI211_X1 g492(.A(new_n689), .B(new_n382), .C1(new_n542), .C2(new_n545), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n542), .B2(new_n545), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n545), .B1(new_n689), .B2(new_n382), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  NOR2_X1   g497(.A1(new_n486), .A2(new_n487), .ZN(new_n699));
  AOI21_X1  g498(.A(G15gat), .B1(new_n689), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n501), .A2(G15gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n689), .B2(new_n701), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n689), .A2(new_n422), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n527), .A2(new_n530), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT84), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT81), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT81), .B1(new_n387), .B2(new_n388), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n422), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n441), .A2(new_n445), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n433), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT78), .B1(new_n520), .B2(new_n521), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n502), .B(new_n382), .C1(new_n519), .C2(new_n428), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n422), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n489), .A2(new_n500), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n390), .A2(new_n447), .A3(KEYINPUT84), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n714), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n706), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n630), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT44), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n566), .A2(new_n687), .A3(new_n660), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n690), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n531), .A2(new_n631), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n570), .A3(new_n690), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT98), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(KEYINPUT45), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(KEYINPUT45), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n571), .A3(new_n382), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT99), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n725), .B2(new_n521), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(G1329gat));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n501), .A3(new_n724), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT100), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n723), .A2(KEYINPUT100), .A3(new_n501), .A4(new_n724), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(G43gat), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n699), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n729), .A2(G43gat), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n742), .B2(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(KEYINPUT47), .B2(new_n751), .ZN(G1330gat));
  NAND3_X1  g551(.A1(new_n723), .A2(new_n422), .A3(new_n724), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n723), .A2(new_n755), .A3(new_n422), .A4(new_n724), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(G50gat), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n711), .A2(G50gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n730), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(KEYINPUT48), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT102), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n753), .A2(new_n764), .A3(G50gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n753), .B2(G50gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n762), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT101), .B(KEYINPUT48), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(G1331gat));
  NOR2_X1   g569(.A1(new_n632), .A2(new_n659), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n721), .A2(new_n687), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n690), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n772), .B(new_n382), .C1(new_n775), .C2(new_n361), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n361), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1333gat));
  XOR2_X1   g577(.A(new_n699), .B(KEYINPUT105), .Z(new_n779));
  AOI21_X1  g578(.A(G71gat), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n718), .A2(new_n480), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n772), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g582(.A1(new_n772), .A2(new_n422), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n726), .A2(G85gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT107), .B1(new_n721), .B2(new_n630), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n789), .B(new_n631), .C1(new_n706), .C2(new_n720), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n566), .A2(new_n659), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT106), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n531), .B2(new_n631), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n721), .A2(KEYINPUT107), .A3(new_n630), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n795), .A2(KEYINPUT51), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT108), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n793), .A3(new_n796), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT108), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n787), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n797), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(KEYINPUT109), .A3(new_n802), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n687), .B(new_n786), .C1(new_n804), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n723), .A2(new_n687), .A3(new_n793), .ZN(new_n810));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810), .B2(new_n726), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1336gat));
  OAI21_X1  g611(.A(G92gat), .B1(new_n810), .B2(new_n521), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n687), .A2(new_n363), .A3(new_n382), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n806), .B2(new_n797), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n799), .B2(new_n803), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(G1337gat));
  NOR2_X1   g620(.A1(new_n747), .A2(G99gat), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n687), .B(new_n822), .C1(new_n804), .C2(new_n808), .ZN(new_n823));
  OAI21_X1  g622(.A(G99gat), .B1(new_n810), .B2(new_n718), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1338gat));
  NAND4_X1  g624(.A1(new_n723), .A2(new_n687), .A3(new_n422), .A4(new_n793), .ZN(new_n826));
  NAND2_X1  g625(.A1(KEYINPUT110), .A2(G106gat), .ZN(new_n827));
  OR2_X1    g626(.A1(KEYINPUT110), .A2(G106gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n687), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n831), .A2(G106gat), .A3(new_n711), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n806), .B2(new_n797), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n799), .B2(new_n803), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(G1339gat));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839));
  INV_X1    g638(.A(new_n566), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n666), .A2(new_n662), .A3(new_n667), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT54), .B(new_n841), .C1(new_n680), .C2(new_n681), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n675), .B1(new_n668), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(KEYINPUT55), .B1(new_n678), .B2(new_n683), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n844), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT111), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n684), .A2(new_n849), .A3(KEYINPUT111), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n659), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n637), .A2(new_n639), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n638), .B1(new_n641), .B2(new_n634), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n654), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n658), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n687), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n630), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n630), .A2(new_n859), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n684), .A2(new_n849), .A3(new_n851), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n865), .B2(new_n852), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n840), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n632), .A2(new_n687), .A3(new_n659), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n839), .B1(new_n870), .B2(new_n711), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n660), .B1(new_n865), .B2(new_n852), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n858), .B1(new_n684), .B2(new_n686), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n631), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n630), .B(new_n859), .C1(new_n850), .C2(new_n853), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n566), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n839), .B(new_n711), .C1(new_n876), .C2(new_n868), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n726), .A2(new_n382), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n699), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n660), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n874), .A2(new_n875), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n868), .B1(new_n885), .B2(new_n840), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n422), .ZN(new_n887));
  INV_X1    g686(.A(new_n881), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n211), .A3(new_n659), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n891), .ZN(G1340gat));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n212), .A3(new_n687), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n212), .B1(new_n882), .B2(new_n687), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1341gat));
  AOI21_X1  g697(.A(G127gat), .B1(new_n890), .B2(new_n566), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n840), .A2(new_n203), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n882), .B2(new_n900), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n883), .B2(new_n631), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n889), .A2(G134gat), .A3(new_n631), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1343gat));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n886), .B2(new_n711), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n847), .A2(new_n909), .A3(new_n848), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n684), .A3(new_n851), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n849), .A2(KEYINPUT115), .B1(new_n657), .B2(new_n658), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n873), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT116), .B1(new_n913), .B2(new_n630), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT55), .B1(new_n842), .B2(new_n844), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n659), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n910), .A2(new_n684), .A3(new_n851), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n860), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n631), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n875), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n868), .B1(new_n921), .B2(new_n840), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n711), .A2(new_n907), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT117), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n912), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n630), .B1(new_n927), .B2(new_n860), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n866), .B1(new_n928), .B2(new_n919), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n566), .B1(new_n929), .B2(new_n914), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n923), .C1(new_n930), .C2(new_n868), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n726), .A2(new_n382), .A3(new_n501), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT114), .Z(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n659), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n906), .B1(new_n935), .B2(G141gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n711), .B1(new_n867), .B2(new_n869), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n933), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(G141gat), .A3(new_n660), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n935), .B2(G141gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n936), .A2(new_n940), .A3(KEYINPUT58), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  AOI221_X4 g741(.A(new_n939), .B1(new_n906), .B2(new_n942), .C1(new_n935), .C2(G141gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(G1344gat));
  NOR4_X1   g743(.A1(new_n501), .A2(G148gat), .A3(new_n831), .A4(new_n711), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n870), .A2(new_n880), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n932), .A2(new_n934), .ZN(new_n947));
  AOI211_X1 g746(.A(KEYINPUT59), .B(new_n227), .C1(new_n947), .C2(new_n687), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT57), .B1(new_n886), .B2(new_n711), .ZN(new_n950));
  INV_X1    g749(.A(new_n928), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n862), .A2(new_n863), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n566), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n907), .B(new_n422), .C1(new_n953), .C2(new_n868), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n950), .A2(new_n687), .A3(new_n934), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n949), .B1(new_n955), .B2(G148gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n946), .B1(new_n948), .B2(new_n956), .ZN(G1345gat));
  NAND3_X1  g756(.A1(new_n947), .A2(G155gat), .A3(new_n566), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n231), .B1(new_n938), .B2(new_n840), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(G1346gat));
  NAND3_X1  g759(.A1(new_n947), .A2(G162gat), .A3(new_n630), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n232), .B1(new_n938), .B2(new_n631), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n690), .A2(new_n521), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n779), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT112), .B1(new_n886), .B2(new_n422), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n877), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G169gat), .B1(new_n968), .B2(new_n660), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n726), .A2(new_n870), .A3(new_n382), .A4(new_n525), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n886), .A2(new_n690), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n382), .A3(new_n525), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT119), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n659), .A2(new_n304), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(G1348gat));
  NOR3_X1   g777(.A1(new_n968), .A2(new_n305), .A3(new_n831), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n831), .B1(new_n972), .B2(new_n975), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n980), .A2(KEYINPUT120), .A3(G176gat), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT120), .B1(new_n980), .B2(G176gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1349gat));
  INV_X1    g782(.A(new_n965), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n566), .B(new_n984), .C1(new_n871), .C2(new_n878), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n967), .A2(new_n987), .A3(new_n566), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(G183gat), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n566), .A3(new_n310), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n970), .A2(KEYINPUT121), .A3(new_n566), .A4(new_n310), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT60), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT60), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n989), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1350gat));
  AOI21_X1  g798(.A(new_n294), .B1(new_n967), .B2(new_n630), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n630), .A2(new_n294), .ZN(new_n1004));
  OAI22_X1  g803(.A1(new_n1002), .A2(new_n1003), .B1(new_n976), .B2(new_n1004), .ZN(G1351gat));
  OAI21_X1  g804(.A(new_n954), .B1(new_n937), .B2(new_n907), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n690), .A2(new_n501), .A3(new_n521), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n954), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n1008), .A2(new_n659), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(G197gat), .ZN(new_n1012));
  AND4_X1   g811(.A1(new_n382), .A2(new_n973), .A3(new_n422), .A4(new_n718), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1013), .A2(new_n340), .A3(new_n659), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(KEYINPUT124), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1012), .A2(new_n1017), .A3(new_n1014), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1016), .A2(new_n1018), .ZN(G1352gat));
  NAND2_X1  g818(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n1013), .A2(new_n341), .A3(new_n687), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g820(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1022));
  XNOR2_X1  g821(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n1024), .A2(new_n687), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1023), .B1(new_n341), .B2(new_n1025), .ZN(G1353gat));
  INV_X1    g825(.A(G211gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1013), .A2(new_n1027), .A3(new_n566), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n950), .A2(new_n566), .A3(new_n954), .A4(new_n1009), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g831(.A(new_n1032), .B(KEYINPUT126), .ZN(G1354gat));
  AOI21_X1  g832(.A(G218gat), .B1(new_n1013), .B2(new_n630), .ZN(new_n1034));
  AND2_X1   g833(.A1(new_n630), .A2(G218gat), .ZN(new_n1035));
  AOI21_X1  g834(.A(new_n1034), .B1(new_n1024), .B2(new_n1035), .ZN(G1355gat));
endmodule


