//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT66), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT2), .A3(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n189), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT67), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT67), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G116), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n190), .A2(new_n192), .B1(new_n188), .B2(new_n189), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n198), .A3(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n202), .A2(new_n204), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G101), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n206), .A2(new_n209), .A3(new_n218), .A4(new_n210), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(KEYINPUT76), .A3(G101), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n198), .A2(KEYINPUT5), .A3(new_n200), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n196), .A2(new_n224), .A3(G116), .A4(new_n197), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(G113), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n198), .A2(new_n200), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n223), .A2(new_n226), .B1(new_n227), .B2(new_n203), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n205), .A2(G107), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n208), .A2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n214), .A2(new_n222), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n187), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n223), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n204), .A3(new_n232), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n211), .A2(new_n213), .A3(G101), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n195), .A2(new_n201), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n193), .A2(new_n194), .B1(new_n198), .B2(new_n200), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n240), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT79), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n235), .B1(new_n238), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT80), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n254), .A2(KEYINPUT64), .A3(G146), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT64), .B1(new_n254), .B2(G146), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n251), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n250), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n253), .B(new_n265), .C1(new_n255), .C2(new_n256), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G143), .B2(new_n252), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n259), .B1(new_n268), .B2(new_n264), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n263), .B1(G125), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT81), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G224), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n275), .B(new_n277), .Z(new_n278));
  NAND2_X1  g092(.A1(new_n246), .A2(KEYINPUT79), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n233), .A2(new_n237), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n187), .A4(new_n236), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n235), .C1(new_n238), .C2(new_n247), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n249), .A2(new_n278), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n275), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n228), .B(new_n232), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n234), .B(KEYINPUT8), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n287), .A2(new_n288), .B1(new_n233), .B2(new_n234), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n284), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n284), .B2(new_n290), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n299));
  NOR2_X1   g113(.A1(G237), .A2(G953), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(G143), .A3(G214), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G143), .B1(new_n300), .B2(G214), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT17), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n276), .A3(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n254), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n301), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT83), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(KEYINPUT16), .A3(G140), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(KEYINPUT16), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n316), .A2(G146), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(G146), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n304), .A2(new_n320), .A3(new_n305), .A4(new_n310), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n304), .A2(new_n305), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n312), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G113), .B(G122), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(new_n205), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n315), .B(new_n252), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT18), .B(G131), .C1(new_n302), .C2(new_n303), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n308), .A2(new_n301), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n304), .A2(new_n310), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n316), .A2(G146), .ZN(new_n333));
  AND2_X1   g147(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n315), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n315), .B2(new_n335), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n332), .B(new_n333), .C1(G146), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n330), .ZN(new_n339));
  INV_X1    g153(.A(new_n325), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G475), .A2(G902), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT84), .A3(KEYINPUT20), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n346));
  INV_X1    g160(.A(new_n343), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n331), .B2(new_n341), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT20), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n342), .B(new_n352), .C1(new_n351), .C2(new_n347), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n323), .A2(new_n330), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n325), .ZN(new_n356));
  OAI21_X1  g170(.A(G475), .B1(new_n356), .B2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT15), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G478), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n254), .A2(G128), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n254), .B2(G128), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n264), .A2(KEYINPUT86), .A3(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G134), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G134), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n371), .A3(new_n362), .ZN(new_n372));
  XNOR2_X1  g186(.A(G116), .B(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n208), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G122), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G116), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n208), .B1(new_n379), .B2(KEYINPUT14), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n377), .A2(KEYINPUT87), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT87), .B1(new_n377), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n373), .A2(new_n208), .ZN(new_n384));
  INV_X1    g198(.A(new_n372), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n371), .B1(new_n368), .B2(new_n362), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n375), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G217), .A3(new_n276), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G902), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n375), .B(new_n391), .C1(new_n383), .C2(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT88), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n398), .A3(new_n394), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n361), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n276), .A2(G952), .ZN(new_n402));
  INV_X1    g216(.A(G234), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n306), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT21), .B(G898), .Z(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT89), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n394), .B(new_n276), .C1(G234), .C2(G237), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT90), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n399), .A2(new_n361), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n299), .B1(new_n358), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n413), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n400), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(KEYINPUT91), .A3(new_n357), .A4(new_n354), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n253), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n258), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n254), .A2(KEYINPUT64), .A3(G146), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n268), .A2(new_n264), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n266), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n232), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n266), .B2(new_n269), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n428), .A2(new_n429), .B1(new_n232), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n257), .A2(new_n261), .A3(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n222), .A2(new_n432), .A3(new_n434), .A4(new_n242), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G137), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT11), .A3(G134), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n371), .A2(G137), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(G134), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT11), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g258(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n437), .C2(G134), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n440), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n440), .B(new_n309), .C1(new_n444), .C2(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n436), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n438), .A2(new_n439), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n441), .A3(new_n443), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n443), .B1(new_n371), .B2(G137), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT65), .ZN(new_n455));
  AOI211_X1 g269(.A(G131), .B(new_n452), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n309), .B1(new_n457), .B2(new_n440), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n431), .A2(new_n435), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n451), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n276), .A2(G227), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT75), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n436), .A2(KEYINPUT77), .A3(new_n449), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n469));
  INV_X1    g283(.A(new_n428), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n232), .A2(new_n270), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n449), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT12), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n449), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n460), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n469), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n461), .A2(new_n469), .A3(new_n466), .A4(new_n467), .ZN(new_n479));
  AOI211_X1 g293(.A(G469), .B(G902), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n461), .A2(new_n467), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n465), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n466), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(G469), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G469), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(new_n394), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n420), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n298), .A2(new_n419), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n442), .A2(new_n439), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G131), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n270), .A2(new_n448), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n432), .A2(new_n434), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT30), .B(new_n495), .C1(new_n496), .C2(new_n459), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n243), .A2(new_n244), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n262), .B1(new_n447), .B2(new_n448), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n270), .A2(new_n448), .A3(new_n494), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n432), .B(new_n434), .C1(new_n456), .C2(new_n458), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n498), .A3(new_n495), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n300), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G101), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n504), .A2(new_n505), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n501), .A2(new_n502), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n498), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(KEYINPUT28), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n516), .A3(new_n498), .A4(new_n495), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n511), .B(KEYINPUT70), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n512), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n504), .A2(new_n507), .A3(new_n511), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT31), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n492), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n518), .A2(new_n520), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n522), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT69), .B1(new_n522), .B2(KEYINPUT31), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n512), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n504), .A2(new_n507), .ZN(new_n537));
  INV_X1    g351(.A(new_n511), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(KEYINPUT71), .A3(new_n538), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT29), .B1(new_n518), .B2(new_n520), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT72), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n498), .B1(new_n506), .B2(new_n495), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n511), .A2(KEYINPUT29), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n546), .B(new_n547), .C1(new_n515), .C2(new_n517), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n548), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n546), .ZN(new_n550));
  INV_X1    g364(.A(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(new_n434), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n433), .B1(new_n257), .B2(new_n261), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n502), .B1(new_n554), .B2(new_n449), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n516), .B1(new_n555), .B2(new_n498), .ZN(new_n556));
  INV_X1    g370(.A(new_n517), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n550), .B(new_n551), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT72), .A3(new_n394), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G472), .B1(new_n544), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n549), .A3(new_n559), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT73), .A3(G472), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n536), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G119), .A2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n196), .A2(new_n197), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(G128), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT24), .B(G110), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n317), .B2(new_n318), .ZN(new_n573));
  INV_X1    g387(.A(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n575));
  AOI21_X1  g389(.A(G128), .B1(new_n196), .B2(new_n197), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n576), .A2(KEYINPUT23), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G140), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G125), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n313), .A2(G140), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n333), .B1(G146), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n575), .A2(new_n574), .A3(new_n577), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n571), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n579), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n573), .A2(new_n578), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n587), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n394), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n592), .A2(KEYINPUT25), .A3(new_n595), .A4(new_n394), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G217), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(G234), .B2(new_n394), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n592), .A2(new_n595), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT74), .B1(new_n567), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n558), .A2(KEYINPUT72), .A3(new_n394), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT72), .B1(new_n558), .B2(new_n394), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n562), .B(new_n609), .C1(new_n612), .C2(new_n564), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT73), .B1(new_n565), .B2(G472), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n530), .B(new_n535), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT74), .ZN(new_n616));
  INV_X1    g430(.A(new_n607), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n491), .B1(new_n608), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n218), .ZN(G3));
  INV_X1    g434(.A(G478), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n396), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n368), .A2(new_n362), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G134), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n372), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n384), .C1(new_n381), .C2(new_n382), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n375), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n392), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT93), .B1(new_n392), .B2(new_n629), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n626), .B2(new_n375), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT33), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n393), .A2(new_n635), .A3(new_n395), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n637), .B(KEYINPUT33), .C1(new_n630), .C2(new_n632), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n394), .A2(G478), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n622), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n358), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n291), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n283), .A2(new_n281), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n279), .A2(new_n280), .A3(new_n236), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n282), .B1(new_n646), .B2(new_n235), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n275), .B(new_n277), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n290), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT92), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n652), .A3(new_n292), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n284), .A2(KEYINPUT92), .A3(new_n290), .A4(new_n291), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n296), .ZN(new_n655));
  AND4_X1   g469(.A1(new_n412), .A2(new_n643), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n609), .B1(new_n534), .B2(new_n394), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n527), .A2(new_n529), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n489), .A2(new_n607), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n401), .A2(new_n413), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n345), .B(new_n350), .C1(KEYINPUT20), .C2(new_n344), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n665), .A3(new_n357), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n412), .A2(new_n653), .A3(new_n655), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n659), .A3(new_n660), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  NAND2_X1  g484(.A1(new_n579), .A2(new_n588), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT96), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n671), .B(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n600), .A2(new_n602), .B1(new_n605), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n657), .A2(new_n658), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n298), .A2(new_n419), .A3(new_n676), .A4(new_n490), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT97), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  NAND2_X1  g494(.A1(new_n563), .A2(new_n566), .ZN(new_n681));
  INV_X1    g495(.A(new_n536), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n675), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n653), .A2(new_n655), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n405), .B1(new_n409), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n666), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n683), .A2(new_n490), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n686), .B(new_n691), .Z(new_n692));
  OR2_X1    g506(.A1(new_n489), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT40), .Z(new_n694));
  AOI21_X1  g508(.A(new_n520), .B1(new_n550), .B2(new_n507), .ZN(new_n695));
  INV_X1    g509(.A(new_n522), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n394), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n295), .B(KEYINPUT38), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n358), .ZN(new_n702));
  INV_X1    g516(.A(new_n675), .ZN(new_n703));
  INV_X1    g517(.A(new_n664), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n297), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n694), .A2(new_n699), .A3(new_n701), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR2_X1   g521(.A1(new_n642), .A2(new_n686), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n683), .A2(new_n490), .A3(new_n684), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n478), .A2(new_n479), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n394), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n485), .A2(KEYINPUT99), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n711), .B(new_n394), .C1(KEYINPUT99), .C2(new_n485), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n420), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n656), .A2(new_n615), .A3(new_n617), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n667), .A2(new_n615), .A3(new_n617), .A4(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  AND2_X1   g536(.A1(new_n415), .A2(new_n418), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n716), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n615), .A3(new_n684), .A4(new_n703), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND3_X1  g540(.A1(new_n358), .A2(new_n412), .A3(new_n664), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT100), .B(G472), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n534), .B2(new_n394), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n696), .A2(new_n505), .B1(new_n519), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n529), .B1(new_n732), .B2(new_n523), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n727), .A2(new_n730), .A3(new_n607), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n684), .A3(new_n717), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  INV_X1    g550(.A(new_n733), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n527), .A2(G902), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n729), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT101), .B1(new_n739), .B2(new_n675), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n534), .A2(new_n394), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n733), .B1(new_n741), .B2(new_n728), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n703), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n653), .A2(new_n655), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n716), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n708), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n651), .A2(new_n296), .A3(new_n292), .A4(new_n420), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n483), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n476), .A2(KEYINPUT102), .A3(new_n466), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n482), .A2(G469), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n487), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n480), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n615), .A2(new_n617), .A3(new_n758), .A4(new_n708), .ZN(new_n759));
  INV_X1    g573(.A(new_n535), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n563), .B2(new_n566), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n534), .A2(new_n528), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(new_n492), .ZN(new_n764));
  AOI211_X1 g578(.A(KEYINPUT103), .B(KEYINPUT32), .C1(new_n534), .C2(new_n528), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n607), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n642), .A2(new_n750), .A3(new_n686), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n750), .A2(new_n759), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n309), .ZN(G33));
  NAND4_X1  g585(.A1(new_n615), .A2(new_n617), .A3(new_n758), .A4(new_n688), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n482), .B2(new_n483), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n485), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n482), .A2(KEYINPUT45), .A3(new_n753), .A4(new_n754), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n486), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT105), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n778), .B(new_n779), .C1(G469), .C2(new_n712), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT104), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n420), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n692), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n702), .A2(new_n641), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n788), .A2(new_n659), .A3(new_n675), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT106), .B(G137), .Z(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  INV_X1    g612(.A(new_n420), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n781), .B2(new_n783), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n708), .A2(new_n793), .A3(new_n607), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n567), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NAND2_X1  g620(.A1(new_n714), .A2(new_n715), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n807), .A2(new_n751), .A3(new_n404), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(new_n788), .ZN(new_n809));
  INV_X1    g623(.A(new_n767), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT48), .Z(new_n812));
  INV_X1    g626(.A(new_n808), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n699), .A2(new_n607), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n643), .A3(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n788), .A2(new_n607), .A3(new_n404), .A4(new_n739), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n747), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n812), .A2(new_n402), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n297), .A3(new_n700), .A4(new_n717), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT50), .B1(new_n819), .B2(KEYINPUT112), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(KEYINPUT112), .B2(new_n819), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n819), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n809), .B1(new_n744), .B2(new_n740), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n813), .A2(new_n814), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n358), .A3(new_n641), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n807), .B(KEYINPUT107), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n799), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n801), .A2(new_n802), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n816), .A2(new_n793), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT111), .Z(new_n833));
  AOI211_X1 g647(.A(new_n826), .B(new_n828), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n818), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n757), .A2(new_n799), .A3(new_n703), .A4(new_n686), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n702), .A2(new_n704), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n699), .A3(new_n684), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n689), .A2(new_n709), .A3(new_n748), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n567), .A2(new_n746), .A3(new_n675), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n490), .C1(new_n688), .C2(new_n708), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n748), .A4(new_n841), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n491), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n567), .A2(KEYINPUT74), .A3(new_n607), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n702), .A2(new_n664), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n411), .B1(new_n853), .B2(new_n642), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n660), .A2(new_n298), .A3(new_n659), .A4(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n735), .A2(new_n855), .A3(new_n677), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n567), .A2(new_n607), .A3(new_n716), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n656), .B2(new_n667), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n852), .A2(new_n856), .A3(new_n858), .A4(new_n725), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n759), .A2(new_n750), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n767), .A2(new_n769), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n743), .B1(new_n742), .B2(new_n703), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n730), .A2(new_n733), .A3(KEYINPUT101), .A4(new_n675), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n708), .B(new_n758), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n664), .A2(new_n686), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n703), .A3(new_n357), .A4(new_n665), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n489), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n615), .A2(new_n868), .A3(new_n793), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n772), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT109), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n865), .A2(new_n772), .A3(new_n869), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n770), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT109), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n735), .A2(new_n855), .A3(new_n677), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n619), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n718), .A2(new_n721), .A3(new_n725), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n875), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n848), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT110), .B1(new_n881), .B2(KEYINPUT53), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n843), .A2(new_n847), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n859), .A2(new_n871), .A3(KEYINPUT109), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n878), .A2(new_n619), .A3(new_n876), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n875), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(KEYINPUT54), .A3(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n859), .A2(new_n871), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n883), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n894), .B(new_n895), .C1(new_n881), .C2(KEYINPUT53), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n838), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n829), .B(KEYINPUT49), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n787), .A2(new_n297), .A3(new_n799), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n700), .A3(new_n814), .A4(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT108), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(G75));
  OAI21_X1  g717(.A(new_n894), .B1(new_n881), .B2(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n394), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n648), .B1(new_n645), .B2(new_n647), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n284), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n912));
  AND3_X1   g726(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n276), .A2(G952), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(G51));
  NAND2_X1  g731(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT116), .A3(new_n896), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n904), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n486), .B(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n711), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n775), .A2(new_n776), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n906), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n916), .B1(new_n924), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n916), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n904), .A2(G902), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n342), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT119), .B1(new_n931), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n904), .A2(G902), .A3(new_n342), .A4(new_n930), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT120), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n933), .B(new_n934), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n929), .A4(new_n940), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(G60));
  XNOR2_X1  g760(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n897), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n639), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  INV_X1    g766(.A(new_n639), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n949), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n919), .A2(new_n921), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n929), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n897), .B2(new_n949), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n929), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT122), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n905), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n674), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n929), .C1(new_n604), .C2(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G66));
  INV_X1    g782(.A(G224), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n408), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n885), .B2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  OAI22_X1  g786(.A1(new_n645), .A2(new_n647), .B1(G898), .B2(new_n276), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(G69));
  AOI21_X1  g788(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n862), .A2(new_n772), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n786), .B2(new_n795), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n845), .A2(new_n748), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n767), .A2(new_n684), .A3(new_n840), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n786), .A2(new_n979), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n805), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n276), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n497), .A2(new_n503), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n337), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n685), .B2(new_n276), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n975), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n978), .A2(new_n706), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n853), .A2(new_n642), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n793), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n693), .B(new_n993), .C1(new_n608), .C2(new_n618), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n786), .B2(new_n795), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n805), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT124), .Z(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n987), .B1(new_n999), .B2(new_n984), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n989), .A2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g815(.A(new_n987), .B1(new_n988), .B2(new_n975), .C1(new_n999), .C2(new_n984), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(new_n537), .A2(new_n511), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n996), .A2(new_n998), .A3(new_n885), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT127), .ZN(new_n1007));
  XOR2_X1   g821(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1004), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1009), .B1(new_n981), .B2(new_n885), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n504), .A2(new_n507), .A3(new_n538), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n929), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n890), .A2(new_n891), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n541), .A2(new_n542), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1009), .B1(new_n1016), .B2(new_n522), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n1011), .B(new_n1014), .C1(new_n1015), .C2(new_n1017), .ZN(G57));
endmodule


