//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203));
  XOR2_X1   g002(.A(G71gat), .B(G99gat), .Z(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G43gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT28), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT68), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(G183gat), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT69), .A4(KEYINPUT28), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n215), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI211_X1 g033(.A(new_n229), .B(new_n234), .C1(KEYINPUT26), .C2(new_n233), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT23), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT24), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT24), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n216), .A3(new_n228), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n242), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n247), .A2(KEYINPUT65), .A3(new_n248), .A4(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n211), .A2(new_n216), .B1(new_n244), .B2(new_n246), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT25), .A4(new_n230), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n221), .A2(new_n216), .A3(new_n222), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n247), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n236), .B1(new_n255), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  INV_X1    g066(.A(G113gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271));
  INV_X1    g070(.A(G134gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G127gat), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n270), .A2(new_n271), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n275), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n257), .A2(new_n256), .A3(new_n258), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n260), .B2(new_n262), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n285), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n243), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n250), .A2(new_n248), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n252), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n242), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n254), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n276), .A2(new_n279), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n236), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n208), .B1(new_n281), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n203), .B(new_n206), .C1(new_n296), .C2(KEYINPUT33), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n206), .A2(new_n203), .A3(KEYINPUT33), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n296), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n281), .A2(new_n295), .A3(new_n208), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT34), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n302), .B1(new_n299), .B2(new_n297), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n307), .B1(new_n300), .B2(new_n303), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT36), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  AND2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(G155gat), .B2(G162gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(new_n280), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n280), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n327), .B2(new_n337), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n337), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT73), .A3(new_n280), .A4(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n294), .A2(new_n338), .A3(KEYINPUT4), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n327), .A2(new_n276), .A3(new_n279), .A4(new_n337), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n341), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n344), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n358), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n350), .B2(new_n353), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n341), .A3(new_n343), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n342), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n320), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n371), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n366), .A2(new_n320), .A3(new_n371), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n377), .B2(KEYINPUT6), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G197gat), .B(G204gat), .Z(new_n385));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G226gat), .ZN(new_n397));
  INV_X1    g196(.A(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n284), .A2(new_n292), .B1(new_n227), .B2(new_n235), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n265), .A2(new_n399), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n265), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n400), .B1(new_n293), .B2(new_n236), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n383), .B1(new_n408), .B2(new_n394), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n388), .A2(new_n384), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n382), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n396), .A3(new_n403), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n406), .B2(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n381), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(KEYINPUT30), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n414), .A2(new_n415), .A3(new_n418), .A4(new_n381), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n376), .A2(new_n378), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n398), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n338), .B1(new_n425), .B2(new_n346), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n347), .A2(new_n405), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n411), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n427), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT3), .B1(new_n396), .B2(new_n405), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n423), .B(new_n430), .C1(new_n431), .C2(new_n338), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT77), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT76), .ZN(new_n437));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(new_n432), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G22gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n435), .A2(new_n442), .A3(new_n434), .A4(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n319), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT37), .B1(new_n404), .B2(new_n412), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n414), .A2(new_n415), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n382), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT38), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n449), .A2(new_n454), .A3(new_n382), .A4(new_n451), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n453), .A2(new_n416), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n376), .A2(new_n378), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n446), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n339), .A2(new_n341), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT39), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n460), .B2(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n360), .A2(KEYINPUT78), .A3(new_n361), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n364), .B2(new_n341), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT79), .B(KEYINPUT39), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n465), .B2(new_n463), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n469), .A2(KEYINPUT80), .A3(new_n371), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT78), .B1(new_n360), .B2(new_n361), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n464), .B(new_n341), .C1(new_n354), .C2(new_n359), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n474), .B2(new_n370), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT40), .B(new_n466), .C1(new_n470), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n466), .B1(new_n470), .B2(new_n475), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT80), .B1(new_n469), .B2(new_n371), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n471), .A3(new_n370), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT40), .A4(new_n466), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n417), .A2(new_n373), .A3(new_n419), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n480), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n458), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n458), .A2(new_n487), .A3(KEYINPUT83), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n448), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n446), .A2(new_n312), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT35), .B1(new_n308), .B2(new_n307), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n421), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n311), .A2(new_n493), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n421), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n311), .A2(new_n493), .A3(KEYINPUT84), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n496), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n202), .B1(new_n492), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n458), .A2(new_n487), .A3(KEYINPUT83), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT83), .B1(new_n458), .B2(new_n487), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n447), .B(new_n319), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n496), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n311), .A2(new_n493), .A3(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT84), .B1(new_n311), .B2(new_n493), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n509), .A2(new_n510), .A3(new_n421), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G43gat), .B(G50gat), .Z(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n524), .B2(KEYINPUT86), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT87), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n518), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n516), .A2(new_n517), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(KEYINPUT87), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n533), .A2(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT17), .A3(new_n529), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G1gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G1gat), .B2(new_n539), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n537), .B2(new_n529), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n544), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT89), .B1(new_n534), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n553), .A2(new_n547), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n546), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n547), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n548), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT12), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n557), .A3(new_n566), .A4(new_n558), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G71gat), .B(G78gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n274), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n544), .B1(new_n574), .B2(new_n573), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT90), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n578), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G155gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n581), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT93), .B(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT8), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(KEYINPUT94), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n600), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n596), .B2(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n602), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n536), .A2(new_n608), .A3(new_n538), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT91), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT41), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n604), .A2(new_n607), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n534), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n612), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT92), .Z(new_n617));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n609), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n609), .B2(new_n615), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n588), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  INV_X1    g423(.A(new_n588), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n620), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n627), .B1(new_n623), .B2(new_n626), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n587), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(G230gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n398), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n603), .B1(new_n636), .B2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g436(.A(new_n573), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n603), .B2(KEYINPUT98), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n606), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n604), .B2(new_n607), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n635), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n638), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n634), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n642), .A2(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n634), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  INV_X1    g453(.A(new_n649), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n646), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT99), .B(new_n654), .C1(new_n646), .C2(new_n655), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n515), .A2(new_n568), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n457), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT100), .B(G1gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1324gat));
  INV_X1    g464(.A(new_n420), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  AND3_X1   g466(.A1(new_n662), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n543), .B1(new_n662), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g470(.A(new_n662), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n672), .A2(G15gat), .A3(new_n316), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n672), .B2(new_n319), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(G1326gat));
  AND2_X1   g474(.A1(new_n515), .A2(new_n568), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n676), .A2(new_n446), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n661), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n631), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n504), .A2(new_n514), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n503), .A2(KEYINPUT103), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n684), .B(new_n496), .C1(new_n502), .C2(KEYINPUT35), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n507), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n629), .A2(new_n630), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n623), .A2(new_n626), .ZN(new_n689));
  INV_X1    g488(.A(new_n627), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT104), .B1(new_n691), .B2(new_n628), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n682), .A2(KEYINPUT44), .B1(new_n686), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n660), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n568), .A3(new_n586), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT102), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n457), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n587), .A2(new_n660), .A3(new_n631), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n515), .A2(new_n568), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n700), .A2(G29gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n704), .A2(new_n702), .A3(new_n706), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n707), .A3(new_n708), .ZN(G1328gat));
  OAI21_X1  g508(.A(G36gat), .B1(new_n699), .B2(new_n420), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n676), .A2(new_n520), .A3(new_n666), .A4(new_n703), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n710), .B(new_n714), .C1(new_n712), .C2(new_n711), .ZN(G1329gat));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n698), .ZN(new_n716));
  INV_X1    g515(.A(new_n319), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(G43gat), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n704), .B2(new_n316), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(new_n446), .ZN(new_n726));
  OAI21_X1  g525(.A(G50gat), .B1(new_n699), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n703), .A2(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n676), .A2(new_n446), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(KEYINPUT48), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n728), .B1(new_n716), .B2(new_n446), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n730), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(G1331gat));
  NOR3_X1   g535(.A1(new_n632), .A2(new_n568), .A3(new_n696), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n686), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n457), .B(KEYINPUT106), .Z(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g542(.A1(new_n738), .A2(new_n420), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  AND2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n744), .B2(new_n745), .ZN(G1333gat));
  NAND3_X1  g547(.A1(new_n739), .A2(G71gat), .A3(new_n717), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n316), .B(KEYINPUT107), .Z(new_n750));
  NOR2_X1   g549(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(G71gat), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n726), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G78gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n587), .A2(new_n631), .A3(new_n568), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT51), .B1(new_n686), .B2(new_n757), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n457), .A3(new_n589), .A4(new_n660), .ZN(new_n761));
  INV_X1    g560(.A(new_n568), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n660), .A2(new_n762), .A3(new_n586), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n695), .A2(new_n700), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  INV_X1    g564(.A(new_n589), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n764), .B2(KEYINPUT109), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n765), .B2(new_n767), .ZN(G1336gat));
  NOR3_X1   g567(.A1(new_n696), .A2(G92gat), .A3(new_n420), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n686), .B2(new_n757), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n758), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(KEYINPUT111), .B(new_n769), .C1(new_n758), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n686), .A2(new_n694), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n763), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n590), .B1(new_n779), .B2(new_n666), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT52), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(new_n760), .B2(new_n769), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(new_n316), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(G99gat), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n760), .A2(new_n786), .A3(new_n660), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n695), .A2(new_n319), .A3(new_n763), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(G1338gat));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n779), .B2(new_n446), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n758), .A2(new_n771), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n696), .A2(G106gat), .A3(new_n726), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT113), .Z(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n779), .B2(new_n446), .ZN(new_n799));
  NOR4_X1   g598(.A1(new_n695), .A2(KEYINPUT114), .A3(new_n726), .A4(new_n763), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n791), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n760), .A2(new_n794), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n801), .B2(new_n804), .ZN(G1339gat));
  NAND2_X1  g604(.A1(new_n568), .A2(new_n268), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT119), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n563), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n567), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n658), .A3(new_n659), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n644), .A2(new_n634), .A3(new_n645), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n815));
  AOI21_X1  g614(.A(new_n652), .B1(new_n646), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n568), .A2(new_n817), .A3(new_n653), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n814), .B2(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n693), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n817), .A2(new_n653), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n814), .A2(new_n816), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n811), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n693), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n586), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n632), .A2(new_n568), .A3(new_n660), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n509), .A2(new_n510), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n741), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT117), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(KEYINPUT118), .A3(new_n420), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT118), .B1(new_n834), .B2(new_n420), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n807), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n700), .A2(new_n666), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n831), .B2(new_n726), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n687), .B1(new_n629), .B2(new_n630), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n691), .A2(KEYINPUT104), .A3(new_n628), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n811), .A3(new_n825), .A4(new_n822), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n693), .A2(new_n820), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n587), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n839), .B(new_n726), .C1(new_n846), .C2(new_n829), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n786), .B(new_n838), .C1(new_n840), .C2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n762), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n837), .A2(new_n850), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n660), .A2(new_n266), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT120), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n835), .B2(new_n836), .ZN(new_n854));
  OAI21_X1  g653(.A(G120gat), .B1(new_n849), .B2(new_n696), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  NAND4_X1  g655(.A1(new_n834), .A2(new_n274), .A3(new_n420), .A4(new_n587), .ZN(new_n857));
  OAI21_X1  g656(.A(G127gat), .B1(new_n849), .B2(new_n586), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  NAND4_X1  g658(.A1(new_n834), .A2(new_n272), .A3(new_n420), .A4(new_n681), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n849), .B2(new_n631), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NOR3_X1   g663(.A1(new_n717), .A2(new_n666), .A3(new_n726), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n831), .A2(new_n741), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n328), .A3(new_n568), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n831), .B2(new_n446), .ZN(new_n869));
  INV_X1    g668(.A(new_n823), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n871));
  OAI211_X1 g670(.A(new_n822), .B(new_n568), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n681), .B1(new_n872), .B2(new_n812), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n586), .B1(new_n873), .B2(new_n827), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n830), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n726), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n869), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n319), .A2(new_n838), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n878), .A2(new_n762), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n868), .B1(new_n880), .B2(new_n328), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n868), .C1(new_n880), .C2(new_n328), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n330), .A3(new_n660), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n878), .A2(new_n696), .A3(new_n879), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(KEYINPUT59), .A3(new_n330), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n826), .A2(new_n631), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n586), .B1(new_n873), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n726), .B1(new_n891), .B2(new_n830), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n844), .A2(new_n845), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n829), .B1(new_n893), .B2(new_n586), .ZN(new_n894));
  INV_X1    g693(.A(new_n877), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n892), .A2(KEYINPUT57), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n696), .B1(new_n879), .B2(KEYINPUT122), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(new_n897), .C1(KEYINPUT122), .C2(new_n879), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n889), .B1(new_n898), .B2(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n886), .B1(new_n888), .B2(new_n899), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n867), .A2(new_n334), .A3(new_n587), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n878), .A2(new_n586), .A3(new_n879), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n334), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n335), .A3(new_n681), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n878), .A2(new_n693), .A3(new_n879), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n335), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n894), .A2(new_n457), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n832), .A2(new_n666), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n568), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n740), .A2(new_n666), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n750), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT116), .B1(new_n894), .B2(new_n446), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n847), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n762), .A2(new_n237), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  NAND3_X1  g718(.A1(new_n911), .A2(new_n238), .A3(new_n660), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n917), .A2(new_n660), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n238), .ZN(G1349gat));
  AND2_X1   g721(.A1(new_n917), .A2(new_n587), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n216), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n587), .A2(new_n212), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  OAI221_X1 g727(.A(new_n928), .B1(new_n910), .B2(new_n925), .C1(new_n923), .C2(new_n216), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n211), .A3(new_n843), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT61), .B(new_n228), .C1(new_n917), .C2(new_n681), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n681), .B(new_n914), .C1(new_n840), .C2(new_n848), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(G190gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n938), .B(new_n931), .C1(new_n932), .C2(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1351gat));
  NAND4_X1  g739(.A1(new_n907), .A2(new_n666), .A3(new_n446), .A4(new_n319), .ZN(new_n941));
  XOR2_X1   g740(.A(KEYINPUT125), .B(G197gat), .Z(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n941), .A2(new_n762), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT126), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n913), .A2(new_n717), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n896), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(new_n762), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(new_n941), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(G204gat), .B1(new_n951), .B2(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n660), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n947), .B2(new_n696), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1353gat));
  OR3_X1    g756(.A1(new_n941), .A2(G211gat), .A3(new_n586), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n896), .A2(new_n587), .A3(new_n946), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n947), .B2(new_n631), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n693), .A2(G218gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n941), .B2(new_n964), .ZN(G1355gat));
endmodule


