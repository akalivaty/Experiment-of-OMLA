//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT69), .Z(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT70), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n464), .A2(G125), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  MUX2_X1   g054(.A(G100), .B(G112), .S(G2105), .Z(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT73), .Z(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n461), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT72), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n482), .A2(new_n488), .A3(new_n493), .ZN(G162));
  NAND2_X1  g069(.A1(new_n492), .A2(G126), .ZN(new_n495));
  MUX2_X1   g070(.A(G102), .B(G114), .S(G2105), .Z(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2104), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n465), .C1(new_n489), .C2(new_n490), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT76), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n486), .A2(new_n502), .A3(new_n503), .A4(G138), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(KEYINPUT74), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n464), .A2(new_n507), .A3(G138), .A4(new_n465), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(KEYINPUT75), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n486), .B2(G138), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n500), .A2(KEYINPUT74), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT4), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n499), .B1(new_n510), .B2(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT77), .Z(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT6), .B(G651), .Z(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n523), .A2(KEYINPUT78), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n529), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n517), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n533), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AND2_X1   g115(.A1(new_n532), .A2(G52), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT79), .B(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n519), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n519), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n532), .A2(G43), .B1(G81), .B2(new_n542), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n532), .A2(new_n562), .A3(G53), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n562), .B1(new_n532), .B2(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT82), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n566), .A2(KEYINPUT83), .A3(new_n519), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT83), .B1(new_n566), .B2(new_n519), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(new_n568), .B1(G91), .B2(new_n542), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n564), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n532), .A2(new_n562), .A3(G53), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  NAND2_X1  g151(.A1(new_n532), .A2(G49), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n517), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n542), .A2(G87), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n517), .A2(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n519), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n542), .A2(G86), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n529), .A2(G48), .A3(G543), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n584), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n519), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT86), .Z(new_n592));
  AOI22_X1  g167(.A1(new_n532), .A2(G47), .B1(G85), .B2(new_n542), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n542), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n532), .A2(G54), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n519), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(G301), .B(new_n601), .S(new_n602), .Z(G284));
  MUX2_X1   g178(.A(G301), .B(new_n601), .S(new_n602), .Z(G321));
  MUX2_X1   g179(.A(G286), .B(G299), .S(new_n602), .Z(G297));
  MUX2_X1   g180(.A(G286), .B(G299), .S(new_n602), .Z(G280));
  AND3_X1   g181(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n601), .A2(G559), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n554), .A2(new_n602), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT11), .Z(G282));
  INV_X1    g189(.A(new_n613), .ZN(G323));
  OAI21_X1  g190(.A(KEYINPUT12), .B1(new_n466), .B2(new_n461), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n486), .A2(new_n617), .A3(G2104), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  MUX2_X1   g198(.A(G99), .B(G111), .S(G2105), .Z(new_n624));
  AOI22_X1  g199(.A1(new_n492), .A2(G123), .B1(G2104), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n466), .ZN(new_n627));
  INV_X1    g202(.A(G2096), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT88), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT89), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  INV_X1    g232(.A(new_n650), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n651), .B(KEYINPUT17), .Z(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n658), .A3(new_n653), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n650), .A3(new_n651), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n628), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n672), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(G166), .A2(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G16), .B2(G22), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT95), .B(G1971), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT94), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n693), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(G6), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G305), .B2(new_n695), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT93), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT32), .B(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G25), .A2(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n492), .A2(G119), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n486), .A2(G131), .ZN(new_n712));
  MUX2_X1   g287(.A(G95), .B(G107), .S(G2105), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2104), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(G16), .A2(G24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G290), .B2(new_n695), .ZN(new_n721));
  INV_X1    g296(.A(G1986), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(new_n721), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n708), .B1(new_n702), .B2(new_n707), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT36), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n726), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n728), .A2(new_n729), .A3(new_n709), .A4(new_n724), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G171), .A2(new_n695), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G5), .B2(new_n695), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n492), .A2(G129), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n486), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n737), .B(new_n740), .C1(G105), .C2(new_n462), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n735), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G34), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n478), .B2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n746), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT100), .Z(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2090), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G2078), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(G16), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n554), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1341), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n757), .A2(new_n760), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n695), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n695), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n695), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n742), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n627), .B2(new_n742), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n744), .B2(new_n745), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n773), .B(new_n778), .C1(new_n734), .C2(new_n733), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n751), .A2(new_n747), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n491), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n465), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n462), .A2(G103), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT25), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT25), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G139), .B2(new_n486), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G33), .B(new_n791), .S(G29), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G2072), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n742), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT28), .Z(new_n795));
  MUX2_X1   g370(.A(G104), .B(G116), .S(G2105), .Z(new_n796));
  AOI22_X1  g371(.A1(new_n492), .A2(G128), .B1(G2104), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n486), .A2(G140), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G4), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n607), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT96), .B(G1348), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n779), .A2(new_n780), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n753), .A2(new_n765), .A3(new_n769), .A4(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n731), .A2(new_n810), .A3(KEYINPUT101), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT101), .B1(new_n731), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(G311));
  NAND2_X1  g388(.A1(new_n731), .A2(new_n810), .ZN(G150));
  NAND2_X1  g389(.A1(new_n532), .A2(G55), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n542), .A2(G93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n815), .B(new_n816), .C1(new_n519), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  OR2_X1    g395(.A1(new_n553), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n553), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n601), .A2(new_n608), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n829), .B2(new_n831), .ZN(G145));
  OAI211_X1 g407(.A(KEYINPUT75), .B(KEYINPUT4), .C1(new_n511), .C2(new_n512), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n501), .A2(new_n504), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n498), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n801), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n715), .B(new_n619), .ZN(new_n839));
  MUX2_X1   g414(.A(G106), .B(G118), .S(G2105), .Z(new_n840));
  AOI22_X1  g415(.A1(new_n492), .A2(G130), .B1(G2104), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G142), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n466), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n838), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n741), .B(new_n791), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n478), .B(new_n627), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n848), .A2(KEYINPUT103), .A3(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n847), .B2(new_n850), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(G395));
  NOR2_X1   g433(.A1(new_n818), .A2(G868), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n823), .A2(new_n610), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n607), .A2(new_n608), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n821), .A3(new_n822), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(G299), .A2(new_n601), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n570), .A2(new_n574), .A3(new_n607), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n607), .B1(new_n570), .B2(new_n574), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT41), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n863), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n860), .A2(new_n864), .A3(new_n866), .A4(new_n862), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT42), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n880), .A2(new_n872), .A3(new_n876), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G288), .ZN(new_n884));
  XNOR2_X1  g459(.A(G303), .B(G305), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n888), .A3(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n859), .B1(new_n890), .B2(G868), .ZN(G295));
  AOI21_X1  g466(.A(new_n859), .B1(new_n890), .B2(G868), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  OR2_X1    g468(.A1(G171), .A2(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g469(.A1(G171), .A2(KEYINPUT107), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(G168), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(G171), .A2(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G286), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n823), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(new_n822), .A3(new_n821), .A4(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n864), .A2(new_n866), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n870), .A2(new_n867), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(new_n902), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(new_n886), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n906), .B2(new_n886), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n902), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(new_n886), .C1(new_n903), .C2(new_n902), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n914), .A2(new_n915), .B1(new_n900), .B2(new_n901), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n870), .A2(KEYINPUT108), .A3(new_n867), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n904), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n912), .B(new_n913), .C1(new_n918), .C2(new_n886), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n893), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n919), .B2(KEYINPUT43), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n918), .A2(new_n886), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(new_n909), .A3(KEYINPUT109), .A4(new_n908), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n922), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n927), .B2(new_n893), .ZN(G397));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G164), .B2(G1384), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n470), .A2(G40), .A3(new_n471), .A4(new_n474), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n801), .B(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT112), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n741), .B(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n715), .B(new_n718), .Z(new_n939));
  OAI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n934), .ZN(new_n941));
  NOR2_X1   g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(KEYINPUT111), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(KEYINPUT111), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT113), .Z(new_n948));
  NAND2_X1  g523(.A1(G303), .A2(G8), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT55), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n931), .B(KEYINPUT110), .ZN(new_n952));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n837), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n930), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1971), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n958));
  INV_X1    g533(.A(G2090), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  NOR3_X1   g535(.A1(G164), .A2(new_n960), .A3(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT50), .B1(new_n837), .B2(new_n953), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n959), .B(new_n952), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n957), .B2(new_n963), .ZN(new_n965));
  OAI211_X1 g540(.A(G8), .B(new_n951), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  NOR2_X1   g542(.A1(G164), .A2(G1384), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n952), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n585), .A2(new_n588), .ZN(new_n970));
  OAI21_X1  g545(.A(G1981), .B1(new_n970), .B2(new_n583), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT116), .B(G1981), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(G305), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT49), .B(new_n971), .C1(G305), .C2(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n952), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n697), .A2(G1976), .ZN(new_n979));
  NAND2_X1  g554(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n978), .A2(G8), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n697), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n969), .B2(new_n979), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n977), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n955), .A2(new_n772), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n747), .B(new_n952), .C1(new_n961), .C2(new_n962), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G8), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G286), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n957), .A2(new_n963), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n950), .B1(new_n993), .B2(new_n967), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n966), .A2(new_n987), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT63), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n964), .B2(new_n965), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n950), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n991), .A2(new_n996), .A3(G286), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n966), .A3(new_n1000), .A4(new_n987), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G288), .A2(G1976), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n977), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G305), .A2(new_n972), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT117), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n969), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n966), .B2(new_n986), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT118), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(new_n1010), .C1(new_n966), .C2(new_n986), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n966), .A2(new_n994), .A3(new_n987), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n955), .B2(G2078), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n734), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n955), .A2(new_n1015), .A3(G2078), .ZN(new_n1020));
  AOI21_X1  g595(.A(G301), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n931), .A2(new_n1015), .A3(G2078), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n930), .A2(new_n954), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(G171), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1014), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n967), .B1(new_n988), .B2(new_n989), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G286), .A2(G8), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT120), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n960), .B1(G164), .B2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n953), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n933), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n747), .A2(new_n1035), .B1(new_n955), .B2(new_n772), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT51), .B(new_n1030), .C1(new_n1036), .C2(new_n967), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n990), .A2(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1032), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1019), .A2(G301), .A3(new_n1020), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1024), .A2(G171), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(KEYINPUT54), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1013), .A2(new_n1026), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2067), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n968), .A2(new_n952), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1045), .B(new_n1046), .C1(new_n1035), .C2(G1348), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1996), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n930), .A2(new_n1049), .A3(new_n954), .A4(new_n952), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n837), .A2(new_n953), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n933), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n554), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT59), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1057), .A3(new_n554), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1048), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n574), .A2(new_n565), .A3(KEYINPUT57), .A4(new_n569), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n569), .B1(new_n564), .B2(new_n563), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1956), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1017), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT56), .B(G2072), .Z(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n930), .A2(new_n952), .A3(new_n954), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1065), .B(new_n1070), .C1(new_n1035), .C2(G1956), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1060), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1017), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n601), .B1(new_n1076), .B2(new_n1045), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n601), .B(new_n1045), .C1(new_n1035), .C2(G1348), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT60), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1070), .B1(new_n1035), .B2(G1956), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT61), .A3(new_n1072), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1059), .A2(new_n1074), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1071), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1002), .B(new_n1012), .C1(new_n1043), .C2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1032), .A2(new_n1037), .A3(new_n1089), .A4(new_n1038), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1021), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n966), .A2(new_n994), .A3(new_n987), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1013), .A2(new_n1094), .A3(new_n1090), .A4(new_n1021), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n948), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n934), .A2(new_n942), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT126), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n940), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n940), .A2(new_n1103), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1101), .B(new_n1102), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n716), .A2(new_n718), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n938), .A2(new_n1107), .B1(G2067), .B2(new_n801), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n934), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n941), .B1(new_n936), .B2(new_n741), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT47), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n934), .B(new_n1049), .C1(KEYINPUT123), .C2(KEYINPUT46), .ZN(new_n1114));
  NAND2_X1  g689(.A1(KEYINPUT123), .A2(KEYINPUT46), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1114), .B(new_n1115), .Z(new_n1116));
  AND3_X1   g691(.A1(new_n1112), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1106), .B(new_n1109), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1097), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g696(.A(G319), .ZN(new_n1123));
  NOR2_X1   g697(.A1(G227), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g698(.A1(new_n1124), .A2(new_n648), .A3(new_n688), .ZN(new_n1125));
  XNOR2_X1  g699(.A(new_n1125), .B(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n856), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g701(.A1(new_n927), .A2(new_n1127), .ZN(G308));
  OR2_X1    g702(.A1(new_n927), .A2(new_n1127), .ZN(G225));
endmodule


