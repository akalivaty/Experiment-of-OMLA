

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597;

  AND2_X1 U328 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U330 ( .A(n421), .B(KEYINPUT11), .ZN(n335) );
  XNOR2_X1 U331 ( .A(n385), .B(n384), .ZN(n541) );
  XNOR2_X1 U332 ( .A(n383), .B(KEYINPUT64), .ZN(n384) );
  XNOR2_X1 U333 ( .A(n298), .B(KEYINPUT13), .ZN(n314) );
  XOR2_X1 U334 ( .A(n311), .B(n336), .Z(n588) );
  XNOR2_X1 U335 ( .A(n386), .B(n296), .ZN(n306) );
  XNOR2_X1 U336 ( .A(n305), .B(n304), .ZN(n307) );
  XNOR2_X1 U337 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U338 ( .A(n342), .B(n341), .ZN(n343) );
  NOR2_X1 U339 ( .A1(n508), .A2(n519), .ZN(n502) );
  XOR2_X1 U340 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n296) );
  XOR2_X1 U341 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n297) );
  INV_X1 U342 ( .A(n572), .ZN(n371) );
  INV_X1 U343 ( .A(KEYINPUT33), .ZN(n302) );
  INV_X1 U344 ( .A(n531), .ZN(n423) );
  XNOR2_X1 U345 ( .A(G71GAT), .B(G78GAT), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U347 ( .A(n333), .B(KEYINPUT78), .ZN(n421) );
  XNOR2_X1 U348 ( .A(n425), .B(KEYINPUT65), .ZN(n582) );
  XNOR2_X1 U349 ( .A(n468), .B(n467), .ZN(n543) );
  XNOR2_X1 U350 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U351 ( .A(n473), .B(n472), .ZN(G1349GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT76), .B(G204GAT), .Z(n429) );
  XNOR2_X1 U353 ( .A(n314), .B(n429), .ZN(n300) );
  AND2_X1 U354 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G148GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n301), .B(G57GAT), .ZN(n414) );
  XNOR2_X1 U358 ( .A(n414), .B(KEYINPUT75), .ZN(n303) );
  XOR2_X1 U359 ( .A(G176GAT), .B(G64GAT), .Z(n386) );
  XOR2_X1 U360 ( .A(KEYINPUT77), .B(G92GAT), .Z(n309) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(n310), .ZN(n336) );
  XNOR2_X1 U364 ( .A(n588), .B(KEYINPUT41), .ZN(n560) );
  XNOR2_X1 U365 ( .A(n560), .B(KEYINPUT108), .ZN(n546) );
  INV_X1 U366 ( .A(n588), .ZN(n354) );
  XOR2_X1 U367 ( .A(KEYINPUT81), .B(G211GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G8GAT), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n398) );
  XNOR2_X1 U370 ( .A(n314), .B(n398), .ZN(n327) );
  XOR2_X1 U371 ( .A(G1GAT), .B(G127GAT), .Z(n416) );
  XOR2_X1 U372 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U373 ( .A(n416), .B(n428), .Z(n316) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U376 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n318) );
  XNOR2_X1 U377 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U379 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U380 ( .A(G15GAT), .B(KEYINPUT73), .Z(n358) );
  XOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n322) );
  XNOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT14), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n358), .B(n323), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n565) );
  XOR2_X1 U387 ( .A(G43GAT), .B(G29GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U390 ( .A(n330), .B(KEYINPUT72), .Z(n332) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n368) );
  XOR2_X1 U393 ( .A(G134GAT), .B(G162GAT), .Z(n333) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n344) );
  INV_X1 U396 ( .A(n336), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n340) );
  XNOR2_X1 U400 ( .A(G190GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n339), .B(KEYINPUT79), .ZN(n392) );
  XOR2_X1 U402 ( .A(n340), .B(n392), .Z(n341) );
  XOR2_X1 U403 ( .A(n368), .B(n345), .Z(n569) );
  INV_X1 U404 ( .A(KEYINPUT80), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n569), .B(n346), .ZN(n348) );
  INV_X1 U406 ( .A(n348), .ZN(n476) );
  INV_X1 U407 ( .A(KEYINPUT36), .ZN(n347) );
  NAND2_X1 U408 ( .A1(n476), .A2(n347), .ZN(n350) );
  NAND2_X1 U409 ( .A1(KEYINPUT36), .A2(n348), .ZN(n349) );
  NAND2_X1 U410 ( .A1(n350), .A2(n349), .ZN(n504) );
  NAND2_X1 U411 ( .A1(n565), .A2(n504), .ZN(n352) );
  XOR2_X1 U412 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  NOR2_X1 U414 ( .A1(n354), .A2(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(KEYINPUT116), .ZN(n372) );
  XOR2_X1 U416 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n357) );
  XNOR2_X1 U417 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U419 ( .A(G197GAT), .B(n358), .Z(n360) );
  XOR2_X1 U420 ( .A(G113GAT), .B(G141GAT), .Z(n417) );
  XNOR2_X1 U421 ( .A(G169GAT), .B(n417), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U424 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n370) );
  XOR2_X1 U426 ( .A(KEYINPUT30), .B(G8GAT), .Z(n366) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(G1GAT), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U429 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n583) );
  XOR2_X1 U431 ( .A(KEYINPUT74), .B(n583), .Z(n572) );
  XNOR2_X1 U432 ( .A(KEYINPUT117), .B(n373), .ZN(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n380) );
  XNOR2_X1 U434 ( .A(n565), .B(KEYINPUT112), .ZN(n574) );
  XOR2_X1 U435 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n376) );
  INV_X1 U436 ( .A(n583), .ZN(n374) );
  NAND2_X1 U437 ( .A1(n560), .A2(n374), .ZN(n375) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n377) );
  NOR2_X1 U439 ( .A1(n574), .A2(n377), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n378), .A2(n569), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  NAND2_X1 U442 ( .A1(n382), .A2(n381), .ZN(n385) );
  INV_X1 U443 ( .A(KEYINPUT48), .ZN(n383) );
  XOR2_X1 U444 ( .A(n386), .B(G92GAT), .Z(n391) );
  XOR2_X1 U445 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U448 ( .A(G169GAT), .B(n389), .Z(n462) );
  XNOR2_X1 U449 ( .A(G36GAT), .B(n462), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n396) );
  XOR2_X1 U451 ( .A(n392), .B(G204GAT), .Z(n394) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U454 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n397), .B(KEYINPUT91), .ZN(n438) );
  XNOR2_X1 U457 ( .A(n438), .B(n398), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n484) );
  NOR2_X1 U459 ( .A1(n541), .A2(n484), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n401), .B(n297), .ZN(n424) );
  XNOR2_X1 U461 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n402), .B(KEYINPUT2), .ZN(n439) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G155GAT), .Z(n404) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(KEYINPUT0), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n406) );
  XNOR2_X1 U467 ( .A(KEYINPUT4), .B(KEYINPUT97), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U469 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n410) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U473 ( .A(KEYINPUT5), .B(n411), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U475 ( .A(n415), .B(n414), .Z(n419) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n439), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n492) );
  XNOR2_X1 U480 ( .A(KEYINPUT99), .B(n492), .ZN(n531) );
  NAND2_X1 U481 ( .A1(n424), .A2(n423), .ZN(n425) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n447) );
  XOR2_X1 U485 ( .A(G162GAT), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n443) );
  XOR2_X1 U488 ( .A(KEYINPUT94), .B(G148GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G50GAT), .B(G106GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U491 ( .A(G78GAT), .B(KEYINPUT93), .Z(n435) );
  XNOR2_X1 U492 ( .A(G141GAT), .B(G211GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n485) );
  NAND2_X1 U501 ( .A1(n582), .A2(n485), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n448), .B(KEYINPUT55), .ZN(n469) );
  XOR2_X1 U503 ( .A(G127GAT), .B(G99GAT), .Z(n450) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G113GAT), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U506 ( .A(G134GAT), .B(G190GAT), .Z(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n466) );
  XOR2_X1 U508 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n454) );
  XNOR2_X1 U509 ( .A(G71GAT), .B(G176GAT), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U511 ( .A(G183GAT), .B(KEYINPUT0), .Z(n456) );
  XNOR2_X1 U512 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U514 ( .A(n458), .B(n457), .Z(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT85), .B(G120GAT), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(n468) );
  NAND2_X1 U521 ( .A1(G227GAT), .A2(G233GAT), .ZN(n467) );
  AND2_X2 U522 ( .A1(n469), .A2(n543), .ZN(n577) );
  AND2_X1 U523 ( .A1(n546), .A2(n577), .ZN(n473) );
  XNOR2_X1 U524 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n471) );
  XNOR2_X1 U525 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n470) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n474) );
  XNOR2_X1 U527 ( .A(n474), .B(KEYINPUT104), .ZN(n475) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(n475), .Z(n498) );
  NAND2_X1 U529 ( .A1(n572), .A2(n588), .ZN(n508) );
  INV_X1 U530 ( .A(n476), .ZN(n576) );
  INV_X1 U531 ( .A(n565), .ZN(n592) );
  NOR2_X1 U532 ( .A1(n576), .A2(n592), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT16), .ZN(n496) );
  XOR2_X1 U534 ( .A(KEYINPUT28), .B(KEYINPUT68), .Z(n478) );
  XNOR2_X1 U535 ( .A(n485), .B(n478), .ZN(n537) );
  XOR2_X1 U536 ( .A(n484), .B(KEYINPUT27), .Z(n483) );
  NAND2_X1 U537 ( .A1(n531), .A2(n483), .ZN(n556) );
  NOR2_X1 U538 ( .A1(n537), .A2(n556), .ZN(n542) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(n542), .ZN(n480) );
  INV_X1 U540 ( .A(n543), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n495) );
  NOR2_X1 U542 ( .A1(n543), .A2(n485), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(n481), .Z(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT26), .B(n482), .ZN(n581) );
  NAND2_X1 U545 ( .A1(n581), .A2(n483), .ZN(n491) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT25), .ZN(n489) );
  INV_X1 U547 ( .A(n484), .ZN(n533) );
  NAND2_X1 U548 ( .A1(n533), .A2(n543), .ZN(n486) );
  NAND2_X1 U549 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n505) );
  NAND2_X1 U555 ( .A1(n496), .A2(n505), .ZN(n519) );
  NAND2_X1 U556 ( .A1(n502), .A2(n531), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U558 ( .A1(n533), .A2(n502), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U561 ( .A1(n502), .A2(n543), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n537), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n505), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n506), .A2(n565), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(KEYINPUT37), .ZN(n528) );
  NOR2_X1 U568 ( .A1(n528), .A2(n508), .ZN(n509) );
  XNOR2_X1 U569 ( .A(KEYINPUT38), .B(n509), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n531), .A2(n517), .ZN(n511) );
  XOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NAND2_X1 U573 ( .A1(n517), .A2(n533), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G36GAT), .B(n513), .ZN(G1329GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n515) );
  NAND2_X1 U577 ( .A1(n543), .A2(n517), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n516), .ZN(G1330GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n537), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n583), .A2(n546), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n529), .A2(n519), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n531), .A2(n524), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n533), .A2(n524), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n543), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U592 ( .A1(n524), .A2(n537), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U594 ( .A(G78GAT), .B(n527), .Z(G1335GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT110), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n536), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U601 ( .A1(n536), .A2(n543), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n541), .A2(n544), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n572), .A2(n552), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  AND2_X1 U611 ( .A1(n546), .A2(n552), .ZN(n548) );
  XNOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(n549), .ZN(G1341GAT) );
  NAND2_X1 U615 ( .A1(n574), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n576), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n555), .Z(G1343GAT) );
  NOR2_X1 U622 ( .A1(n541), .A2(n556), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n557), .A2(n581), .ZN(n568) );
  NOR2_X1 U624 ( .A1(n583), .A2(n568), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(n558), .Z(n559) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT121), .Z(n562) );
  INV_X1 U628 ( .A(n568), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  OR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT122), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G162GAT), .B(n571), .ZN(G1347GAT) );
  AND2_X1 U638 ( .A1(n572), .A2(n577), .ZN(n573) );
  XOR2_X1 U639 ( .A(G169GAT), .B(n573), .Z(G1348GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(n580), .ZN(G1351GAT) );
  XNOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n594) );
  NOR2_X1 U648 ( .A1(n583), .A2(n594), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n594), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(G204GAT), .B(n591), .Z(G1353GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n594), .ZN(n593) );
  XOR2_X1 U657 ( .A(G211GAT), .B(n593), .Z(G1354GAT) );
  INV_X1 U658 ( .A(n594), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n504), .A2(n595), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

