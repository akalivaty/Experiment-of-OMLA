

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U325 ( .A(n432), .B(n309), .Z(n537) );
  XNOR2_X1 U326 ( .A(n327), .B(n326), .ZN(n526) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n403) );
  XOR2_X1 U328 ( .A(KEYINPUT111), .B(n412), .Z(n292) );
  INV_X1 U329 ( .A(KEYINPUT88), .ZN(n463) );
  XNOR2_X1 U330 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U331 ( .A1(n465), .A2(n473), .ZN(n467) );
  INV_X1 U332 ( .A(KEYINPUT32), .ZN(n366) );
  XNOR2_X1 U333 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U334 ( .A(n389), .B(n368), .ZN(n369) );
  INV_X1 U335 ( .A(KEYINPUT11), .ZN(n390) );
  NOR2_X1 U336 ( .A1(n563), .A2(n493), .ZN(n494) );
  XNOR2_X1 U337 ( .A(n404), .B(KEYINPUT36), .ZN(n405) );
  XNOR2_X1 U338 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U339 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U340 ( .A(n406), .B(n405), .ZN(n492) );
  XNOR2_X1 U341 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n453) );
  NOR2_X1 U342 ( .A1(n492), .A2(n495), .ZN(n496) );
  XNOR2_X1 U343 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U344 ( .A1(n537), .A2(n455), .ZN(n571) );
  XOR2_X1 U345 ( .A(n434), .B(n433), .Z(n524) );
  XNOR2_X1 U346 ( .A(KEYINPUT38), .B(n498), .ZN(n506) );
  XNOR2_X1 U347 ( .A(n460), .B(G190GAT), .ZN(n461) );
  XOR2_X1 U348 ( .A(G127GAT), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U349 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(n295), .ZN(n432) );
  XOR2_X1 U352 ( .A(G99GAT), .B(G43GAT), .Z(n297) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n300) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n312) );
  XOR2_X1 U358 ( .A(n300), .B(n312), .Z(n308) );
  XOR2_X1 U359 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n302) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U362 ( .A(G183GAT), .B(G71GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(G15GAT), .B(G176GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U367 ( .A(G211GAT), .B(KEYINPUT83), .Z(n311) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n448) );
  XNOR2_X1 U370 ( .A(n312), .B(n448), .ZN(n327) );
  XOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .Z(n331) );
  INV_X1 U372 ( .A(KEYINPUT77), .ZN(n313) );
  NAND2_X1 U373 ( .A1(n313), .A2(G218GAT), .ZN(n316) );
  INV_X1 U374 ( .A(G218GAT), .ZN(n314) );
  NAND2_X1 U375 ( .A1(n314), .A2(KEYINPUT77), .ZN(n315) );
  NAND2_X1 U376 ( .A1(n316), .A2(n315), .ZN(n318) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n392) );
  XOR2_X1 U379 ( .A(KEYINPUT87), .B(n392), .Z(n322) );
  XOR2_X1 U380 ( .A(G64GAT), .B(KEYINPUT73), .Z(n320) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G204GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n373) );
  XNOR2_X1 U383 ( .A(n373), .B(G92GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U385 ( .A(n331), .B(n323), .Z(n325) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U388 ( .A(KEYINPUT109), .B(KEYINPUT47), .Z(n402) );
  XOR2_X1 U389 ( .A(KEYINPUT15), .B(G64GAT), .Z(n329) );
  XNOR2_X1 U390 ( .A(G127GAT), .B(G211GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n344) );
  XNOR2_X1 U392 ( .A(G71GAT), .B(G57GAT), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n330), .B(KEYINPUT13), .ZN(n372) );
  XOR2_X1 U394 ( .A(n372), .B(n331), .Z(n333) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U397 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n335) );
  XNOR2_X1 U398 ( .A(KEYINPUT14), .B(KEYINPUT78), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U400 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U401 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n339) );
  XNOR2_X1 U402 ( .A(G15GAT), .B(G1GAT), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n356) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n340), .B(G78GAT), .ZN(n440) );
  XNOR2_X1 U406 ( .A(n356), .B(n440), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n587) );
  XOR2_X1 U409 ( .A(KEYINPUT106), .B(n587), .Z(n572) );
  XOR2_X1 U410 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n346) );
  XNOR2_X1 U411 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n363) );
  XOR2_X1 U413 ( .A(G113GAT), .B(G36GAT), .Z(n348) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G50GAT), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U416 ( .A(G8GAT), .B(G22GAT), .Z(n350) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G141GAT), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U419 ( .A(n352), .B(n351), .Z(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n354) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G29GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(n355), .Z(n388) );
  XOR2_X1 U424 ( .A(n356), .B(KEYINPUT71), .Z(n358) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n388), .B(n359), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n569) );
  INV_X1 U430 ( .A(n569), .ZN(n577) );
  XOR2_X1 U431 ( .A(KEYINPUT72), .B(G92GAT), .Z(n365) );
  XNOR2_X1 U432 ( .A(G99GAT), .B(G85GAT), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n389) );
  NAND2_X1 U434 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n369), .B(G78GAT), .ZN(n371) );
  XOR2_X1 U436 ( .A(G106GAT), .B(G148GAT), .Z(n437) );
  XOR2_X1 U437 ( .A(G120GAT), .B(n437), .Z(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U440 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n375) );
  XNOR2_X1 U441 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U443 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n403), .B(n380), .ZN(n543) );
  NOR2_X1 U445 ( .A1(n577), .A2(n543), .ZN(n382) );
  XNOR2_X1 U446 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U448 ( .A(KEYINPUT107), .B(n383), .Z(n384) );
  NOR2_X1 U449 ( .A1(n572), .A2(n384), .ZN(n400) );
  XOR2_X1 U450 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n386) );
  XNOR2_X1 U451 ( .A(G134GAT), .B(G106GAT), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U453 ( .A(n388), .B(n387), .Z(n398) );
  XNOR2_X1 U454 ( .A(n389), .B(KEYINPUT76), .ZN(n391) );
  XOR2_X1 U455 ( .A(G50GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U456 ( .A(n392), .B(n439), .ZN(n394) );
  AND2_X1 U457 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n406) );
  INV_X1 U460 ( .A(n406), .ZN(n399) );
  NAND2_X1 U461 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n413) );
  INV_X1 U463 ( .A(KEYINPUT45), .ZN(n408) );
  INV_X1 U464 ( .A(KEYINPUT96), .ZN(n404) );
  NOR2_X1 U465 ( .A1(n492), .A2(n587), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  NOR2_X1 U467 ( .A1(n403), .A2(n409), .ZN(n410) );
  XOR2_X1 U468 ( .A(KEYINPUT110), .B(n410), .Z(n411) );
  NOR2_X1 U469 ( .A1(n569), .A2(n411), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n413), .A2(n292), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(KEYINPUT48), .ZN(n534) );
  NOR2_X1 U472 ( .A1(n526), .A2(n534), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n415), .B(KEYINPUT54), .ZN(n435) );
  XOR2_X1 U474 ( .A(G57GAT), .B(KEYINPUT6), .Z(n417) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n431) );
  XOR2_X1 U477 ( .A(KEYINPUT84), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U478 ( .A(G148GAT), .B(G162GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n421) );
  XNOR2_X1 U481 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n429) );
  XNOR2_X1 U484 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n424), .B(KEYINPUT2), .ZN(n447) );
  XOR2_X1 U486 ( .A(G85GAT), .B(n447), .Z(n426) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n434) );
  INV_X1 U492 ( .A(n432), .ZN(n433) );
  NAND2_X1 U493 ( .A1(n435), .A2(n524), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n436), .B(KEYINPUT65), .ZN(n576) );
  XNOR2_X1 U495 ( .A(G218GAT), .B(G204GAT), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n452) );
  XOR2_X1 U497 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n444) );
  XNOR2_X1 U501 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n473) );
  NAND2_X1 U507 ( .A1(n576), .A2(n473), .ZN(n454) );
  INV_X1 U508 ( .A(n543), .ZN(n558) );
  NAND2_X1 U509 ( .A1(n571), .A2(n558), .ZN(n459) );
  XOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT122), .Z(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  NAND2_X1 U514 ( .A1(n571), .A2(n406), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n460) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  NOR2_X1 U517 ( .A1(n577), .A2(n403), .ZN(n497) );
  NOR2_X1 U518 ( .A1(n526), .A2(n537), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(KEYINPUT89), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n467), .B(n466), .ZN(n470) );
  INV_X1 U521 ( .A(n537), .ZN(n474) );
  NOR2_X1 U522 ( .A1(n473), .A2(n474), .ZN(n468) );
  XOR2_X1 U523 ( .A(n468), .B(KEYINPUT26), .Z(n574) );
  XNOR2_X1 U524 ( .A(n526), .B(KEYINPUT27), .ZN(n533) );
  OR2_X1 U525 ( .A1(n574), .A2(n533), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT90), .B(n471), .Z(n472) );
  NAND2_X1 U528 ( .A1(n472), .A2(n524), .ZN(n478) );
  INV_X1 U529 ( .A(n524), .ZN(n536) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(n473), .ZN(n539) );
  NOR2_X1 U531 ( .A1(n533), .A2(n474), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n539), .A2(n475), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n536), .A2(n476), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n493) );
  NOR2_X1 U535 ( .A1(n406), .A2(n587), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U537 ( .A1(n493), .A2(n480), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT91), .B(n481), .Z(n510) );
  NAND2_X1 U539 ( .A1(n497), .A2(n510), .ZN(n490) );
  NOR2_X1 U540 ( .A1(n524), .A2(n490), .ZN(n482) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n482), .Z(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n526), .A2(n490), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n537), .A2(n490), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n539), .A2(n490), .ZN(n491) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  INV_X1 U553 ( .A(n587), .ZN(n563) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT97), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT37), .B(n496), .Z(n523) );
  NAND2_X1 U556 ( .A1(n523), .A2(n497), .ZN(n498) );
  NOR2_X1 U557 ( .A1(n506), .A2(n524), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT95), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n502) );
  XOR2_X1 U560 ( .A(KEYINPUT39), .B(KEYINPUT98), .Z(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n526), .A2(n506), .ZN(n503) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U564 ( .A1(n506), .A2(n537), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(n504), .Z(n505) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  XNOR2_X1 U567 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n508) );
  NOR2_X1 U568 ( .A1(n539), .A2(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  NOR2_X1 U571 ( .A1(n569), .A2(n543), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n522), .A2(n510), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n524), .A2(n519), .ZN(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT101), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n526), .A2(n519), .ZN(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n537), .A2(n519), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  NOR2_X1 U584 ( .A1(n539), .A2(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n524), .A2(n530), .ZN(n525) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n526), .A2(n530), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n537), .A2(n530), .ZN(n529) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n539), .A2(n530), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n555) );
  NOR2_X1 U600 ( .A1(n537), .A2(n555), .ZN(n538) );
  XNOR2_X1 U601 ( .A(KEYINPUT112), .B(n538), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n577), .A2(n547), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  NOR2_X1 U606 ( .A1(n543), .A2(n547), .ZN(n545) );
  XNOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n549) );
  INV_X1 U611 ( .A(n547), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n551), .A2(n572), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U616 ( .A1(n551), .A2(n406), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT117), .Z(n557) );
  NOR2_X1 U620 ( .A1(n574), .A2(n555), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n565), .A2(n569), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U625 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n567) );
  NAND2_X1 U631 ( .A1(n565), .A2(n406), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n571), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U638 ( .A(n574), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n589) );
  NOR2_X1 U640 ( .A1(n577), .A2(n589), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  INV_X1 U644 ( .A(n403), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n581), .A2(n589), .ZN(n586) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT124), .B(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n589), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n492), .A2(n589), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

