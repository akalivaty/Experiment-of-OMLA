//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT70), .Z(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT71), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(G567), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT73), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G113), .A3(G2104), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n467), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n471), .B1(new_n470), .B2(new_n474), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n468), .A2(new_n469), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(new_n467), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  AND2_X1   g065(.A1(G112), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G100), .B2(new_n467), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n488), .B(new_n490), .C1(new_n472), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT75), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND2_X1  g070(.A1(new_n467), .A2(G102), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n472), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n468), .B2(new_n469), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(KEYINPUT76), .B(new_n499), .C1(new_n468), .C2(new_n469), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT3), .B(G2104), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G138), .A4(new_n467), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(G50), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(new_n513), .B2(new_n514), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(G62), .B1(new_n517), .B2(new_n516), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT77), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n523), .ZN(new_n530));
  OAI21_X1  g105(.A(G651), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(new_n528), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(new_n535), .A3(G88), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n531), .A2(new_n536), .A3(new_n537), .A4(new_n515), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(new_n538), .ZN(G166));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n517), .A2(new_n516), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n534), .A2(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(G63), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n521), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(new_n553), .B2(new_n552), .ZN(new_n555));
  INV_X1    g130(.A(new_n518), .ZN(new_n556));
  INV_X1    g131(.A(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n532), .B2(new_n533), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n556), .A2(G90), .B1(new_n558), .B2(G52), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n521), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n556), .A2(G81), .B1(new_n558), .B2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT79), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n558), .B(G53), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n545), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(G651), .A2(new_n581), .B1(new_n556), .B2(G91), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n525), .A2(new_n585), .A3(new_n538), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n525), .B2(new_n538), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n586), .A2(new_n587), .ZN(G303));
  NAND2_X1  g163(.A1(new_n556), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n558), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n556), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n558), .A2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n535), .A2(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n521), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n521), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n542), .A2(new_n603), .B1(new_n518), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n535), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n521), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n518), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n558), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n558), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g195(.A(G54), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n609), .B1(new_n622), .B2(new_n608), .ZN(G284));
  XNOR2_X1  g198(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NOR2_X1   g199(.A1(G286), .A2(new_n608), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n608), .ZN(G297));
  AOI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(new_n608), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NOR2_X1   g205(.A1(new_n565), .A2(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n616), .A2(new_n621), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G559), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n631), .B1(new_n633), .B2(G868), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n487), .A2(G2104), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT84), .B(G2100), .Z(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  MUX2_X1   g216(.A(G99), .B(G111), .S(G2105), .Z(new_n642));
  AOI22_X1  g217(.A1(new_n489), .A2(G123), .B1(G2104), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n507), .A2(new_n467), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n641), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2427), .ZN(new_n652));
  INV_X1    g227(.A(G2430), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n656), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT86), .Z(new_n665));
  INV_X1    g240(.A(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  INV_X1    g251(.A(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .A3(new_n670), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n670), .B1(new_n677), .B2(KEYINPUT17), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n671), .A2(new_n674), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n681), .B2(KEYINPUT17), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n647), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT89), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  NAND2_X1  g281(.A1(new_n606), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n487), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n489), .A2(G119), .ZN(new_n712));
  MUX2_X1   g287(.A(G95), .B(G107), .S(G2105), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2104), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G25), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT90), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n718), .A2(new_n721), .B1(new_n708), .B2(new_n709), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n710), .B(new_n722), .C1(new_n718), .C2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G22), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT93), .B(G1971), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G6), .A2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n599), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n724), .A2(G23), .ZN(new_n734));
  INV_X1    g309(.A(G288), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n724), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT33), .B(G1976), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n729), .A2(new_n733), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n723), .B1(new_n740), .B2(KEYINPUT34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(KEYINPUT34), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n724), .A2(G20), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT23), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n724), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n724), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1961), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G160), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n753), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n751), .B1(G1961), .B2(new_n749), .C1(new_n752), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n753), .A2(G35), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n494), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT97), .B(G28), .Z(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(KEYINPUT30), .B2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n768), .B(new_n769), .C1(new_n646), .C2(new_n753), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n724), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n724), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(new_n772), .B2(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n622), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G4), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1348), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n773), .B1(G1966), .B2(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n758), .A2(new_n752), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR4_X1    g355(.A1(new_n759), .A2(new_n765), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT96), .B1(G29), .B2(G32), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n487), .A2(G141), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n489), .A2(G129), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G105), .B2(new_n473), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n753), .ZN(new_n795));
  MUX2_X1   g370(.A(new_n783), .B(KEYINPUT96), .S(new_n795), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G19), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n566), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1341), .ZN(new_n802));
  NOR2_X1   g377(.A1(G27), .A2(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G164), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2078), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n753), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n487), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n489), .A2(G128), .ZN(new_n809));
  MUX2_X1   g384(.A(G104), .B(G116), .S(G2105), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2104), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n753), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2067), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n802), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G29), .A2(G33), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT25), .B1(new_n473), .B2(G103), .ZN(new_n820));
  INV_X1    g395(.A(G139), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n819), .A2(new_n820), .B1(new_n645), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n507), .A2(G127), .ZN(new_n823));
  NAND2_X1  g398(.A1(G115), .A2(G2104), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n467), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n817), .B1(new_n826), .B2(G29), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT94), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2072), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n798), .A2(new_n799), .A3(new_n816), .A4(new_n829), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n781), .A2(new_n782), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n782), .B1(new_n781), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n743), .B1(new_n831), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n743), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  AOI22_X1  g411(.A1(new_n556), .A2(G93), .B1(new_n558), .B2(G55), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n521), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n565), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n565), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n622), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n841), .B1(new_n850), .B2(new_n852), .ZN(G145));
  INV_X1    g428(.A(new_n826), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT102), .B1(new_n854), .B2(KEYINPUT101), .ZN(new_n855));
  INV_X1    g430(.A(new_n794), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n813), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n794), .A2(new_n812), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G164), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n511), .A3(new_n858), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n637), .B(new_n715), .ZN(new_n865));
  MUX2_X1   g440(.A(G106), .B(G118), .S(G2105), .Z(new_n866));
  AOI22_X1  g441(.A1(new_n489), .A2(G130), .B1(G2104), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n645), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n865), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n861), .A2(new_n863), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(new_n860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n855), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n494), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n646), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n864), .A2(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n872), .A3(new_n860), .ZN(new_n879));
  INV_X1    g454(.A(new_n855), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n875), .A2(new_n884), .A3(new_n877), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n877), .B1(new_n875), .B2(new_n881), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(G37), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT40), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(G395));
  NAND2_X1  g466(.A1(new_n622), .A2(new_n626), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n632), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n844), .B1(G559), .B2(new_n632), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n842), .A2(new_n843), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n633), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n894), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n896), .A2(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n899), .A2(new_n894), .A3(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G166), .B(new_n599), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n735), .B(new_n606), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n911), .B(new_n912), .Z(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n906), .A2(new_n909), .A3(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(G868), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n920), .A3(G868), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n839), .A2(new_n608), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n608), .B1(new_n910), .B2(new_n915), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n925), .B2(new_n917), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT106), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n919), .A2(new_n928), .A3(new_n921), .A4(new_n922), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g506(.A(G301), .B(G168), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(new_n844), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n844), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n933), .A2(new_n934), .A3(new_n894), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n896), .B(new_n897), .C1(new_n933), .C2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT108), .A3(new_n913), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n913), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n941), .A3(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n913), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n931), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n939), .A3(new_n942), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT44), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT107), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n940), .A2(new_n945), .A3(new_n931), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n949), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n511), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n481), .A2(new_n482), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G2105), .ZN(new_n963));
  INV_X1    g538(.A(new_n484), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(G40), .A4(new_n475), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G2067), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n812), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n856), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT46), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n856), .A2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n794), .A2(G1996), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n969), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n716), .A2(new_n719), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(G2067), .B2(new_n812), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n966), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n966), .A2(new_n709), .A3(new_n606), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  INV_X1    g559(.A(new_n979), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n716), .A2(new_n719), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n980), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n988), .B2(new_n967), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n976), .A2(new_n982), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n965), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n504), .B2(new_n510), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n961), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT56), .B(G2072), .Z(new_n995));
  OR2_X1    g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n997));
  NAND2_X1  g572(.A1(G299), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n578), .A2(KEYINPUT121), .A3(new_n999), .A4(new_n582), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n992), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(G160), .B(G40), .C1(new_n992), .C2(new_n1004), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1003), .B1(new_n992), .B2(new_n1004), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n996), .B(new_n1002), .C1(G1956), .C2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT50), .B(G1384), .C1(new_n504), .C2(new_n510), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n776), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n959), .A2(new_n965), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n968), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n632), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n965), .B1(new_n959), .B2(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1956), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n994), .A2(new_n995), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1001), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT58), .B(G1341), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(G160), .B(G40), .C1(new_n992), .C2(KEYINPUT45), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1027), .B2(new_n972), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT59), .B1(new_n1028), .B2(new_n565), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n994), .A2(G1996), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1030), .B(new_n566), .C1(new_n1031), .C2(new_n1024), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1012), .A2(new_n632), .A3(new_n1014), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT60), .B1(new_n1034), .B2(new_n1015), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n632), .A2(KEYINPUT60), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1012), .A2(new_n1036), .A3(new_n1014), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT61), .B1(new_n1021), .B2(new_n1010), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1021), .A2(new_n1010), .A3(KEYINPUT61), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT122), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1021), .A2(new_n1010), .A3(new_n1043), .A4(KEYINPUT61), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1022), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(KEYINPUT109), .B2(KEYINPUT55), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n586), .B2(new_n587), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g628(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .C1(new_n586), .C2(new_n587), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n511), .A2(new_n1004), .A3(new_n958), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1018), .A2(new_n1058), .A3(new_n764), .A4(new_n1005), .ZN(new_n1059));
  INV_X1    g634(.A(G1971), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1056), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT117), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1064), .A2(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n965), .B1(new_n959), .B2(new_n960), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1971), .B1(new_n1068), .B2(new_n993), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1007), .A2(G2090), .A3(new_n1011), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1018), .A2(new_n764), .A3(new_n1057), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1056), .B1(new_n1061), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT110), .B1(new_n1055), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1063), .B(new_n1067), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n735), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n991), .A2(new_n992), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n959), .B2(new_n965), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1081), .A2(new_n1084), .B1(G1976), .B2(new_n735), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(KEYINPUT112), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1079), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n735), .A2(G1976), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1087), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n598), .ZN(new_n1095));
  INV_X1    g670(.A(G1981), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n593), .A4(new_n594), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT113), .B(G86), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n594), .B1(new_n518), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1099), .B2(new_n598), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n1100), .A3(KEYINPUT49), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT49), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT111), .B1(new_n1080), .B2(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n1103), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1094), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1078), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n1113));
  INV_X1    g688(.A(G1966), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n994), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1018), .A2(new_n1116), .A3(new_n752), .A4(new_n1057), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1119), .B2(new_n752), .ZN(new_n1120));
  OAI21_X1  g695(.A(G8), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G168), .A2(new_n1056), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n1123), .B2(KEYINPUT123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1018), .A2(new_n1057), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT118), .B1(new_n1127), .B2(G2084), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(new_n1117), .A3(new_n1115), .ZN(new_n1129));
  OAI211_X1 g704(.A(G8), .B(new_n1124), .C1(new_n1129), .C2(G286), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(G8), .A3(G286), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G301), .B(KEYINPUT54), .ZN(new_n1133));
  INV_X1    g708(.A(G2078), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1134), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n964), .A2(new_n475), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n962), .B(KEYINPUT125), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(G2105), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(new_n961), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1133), .B1(new_n993), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1068), .A2(new_n1134), .A3(new_n993), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  INV_X1    g717(.A(G1961), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1141), .A2(new_n1142), .B1(new_n1127), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT53), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1144), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1149), .B2(new_n1133), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1112), .A2(new_n1113), .A3(new_n1132), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1132), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1073), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1076), .A2(KEYINPUT110), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1153), .A2(new_n1154), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1088), .A2(new_n1093), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1063), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT126), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1046), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1076), .A2(KEYINPUT120), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1076), .A2(KEYINPUT120), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1072), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1121), .A2(G286), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT63), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1164), .A2(new_n1166), .A3(new_n1111), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1155), .A2(new_n1156), .A3(new_n1163), .A4(new_n1063), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n1168), .B2(KEYINPUT119), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1078), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1156), .A4(new_n1163), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1132), .A2(KEYINPUT62), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1126), .A2(new_n1130), .A3(new_n1175), .A4(new_n1131), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1148), .B2(new_n1144), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1112), .A2(new_n1174), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1111), .A2(new_n1165), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1089), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1097), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1110), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1180), .B1(new_n1183), .B2(KEYINPUT115), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT115), .ZN(new_n1185));
  AOI211_X1 g760(.A(G1976), .B(G288), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n1181), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1179), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1178), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1159), .A2(new_n1173), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n606), .B(G1986), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n967), .B1(new_n988), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n990), .B1(new_n1190), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g768(.A1(new_n886), .A2(new_n888), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n465), .A2(G227), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n668), .A2(new_n705), .A3(new_n1197), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(G308));
  NAND3_X1  g773(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(G225));
endmodule


